// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

         if(local_pf_num == 'h0 && local_vf_num == 'd0 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D0, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;
                                                                                              })

        `reset_in_middle(0)

 	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd3 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D3, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(3)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd4 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D4, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(4)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd5 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D5, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(5)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd6 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D6, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(6)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd7 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D7, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(7)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd8 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D8, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(8)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd9 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D9, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(9)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd10 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D10, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(10)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd11 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D11, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(11)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd12 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D12, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(12)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd13 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D13, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(13)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd14 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D14, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(14)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd15 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D15, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(15)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd16 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D16, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(16)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd17 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D17, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(17)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd18 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D18, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(18)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd19 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D19, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(19)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd20 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D20, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(20)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd21 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D21, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(21)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd22 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D22, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(22)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd23 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D23, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(23)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd24 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D24, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(24)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd25 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D25, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(25)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd26 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D26, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(26)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd27 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D27, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(27)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd28 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D28, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(28)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd29 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D29, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(29)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd30 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D30, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(30)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd31 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D31, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(31)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd32 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D32, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(32)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd33 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D33, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(33)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd34 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D34, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(34)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd35 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D35, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(35)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd36 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D36, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(36)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd37 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D37, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(37)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd38 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D38, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(38)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd39 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D39, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(39)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd40 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D40, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(40)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd41 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D41, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(41)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd42 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D42, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(42)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd43 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D43, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(43)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd44 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D44, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(44)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd45 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D45, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(45)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd46 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D46, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(46)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd47 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D47, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(47)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd48 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D48, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(48)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd49 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D49, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(49)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd50 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D50, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(50)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd51 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D51, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(51)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd52 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D52, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(52)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd53 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D53, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(53)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd54 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D54, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(54)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd55 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D55, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(55)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd56 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D56, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(56)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd57 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D57, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(57)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd58 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D58, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(58)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd59 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D59, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(59)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd60 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D60, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(60)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd61 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D61, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(61)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd62 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D62, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(62)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd63 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D63, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(63)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd64 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D64, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(64)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd65 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D65, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(65)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd66 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D66, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(66)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd67 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D67, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(67)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd68 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D68, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(68)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd69 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D69, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(69)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd70 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D70, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(70)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd71 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D71, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(71)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd72 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D72, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(72)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd73 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D73, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(73)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd74 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D74, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(74)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd75 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D75, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(75)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd76 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D76, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(76)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd77 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D77, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(77)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd78 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D78, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(78)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd79 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D79, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(79)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd80 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D80, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(80)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd81 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D81, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(81)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd82 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D82, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(82)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd83 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D83, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(83)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd84 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D84, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(84)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd85 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D85, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(85)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd86 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D86, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(86)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd87 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D87, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(87)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd88 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D88, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(88)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd89 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D89, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(89)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd90 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D90, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(90)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd91 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D91, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(91)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd92 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D92, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(92)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd93 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D93, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(93)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd94 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D94, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(94)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd95 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D95, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(95)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd96 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D96, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(96)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd97 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D97, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(97)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd98 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D98, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(98)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd99 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D99, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(99)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd100 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(100)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd101 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(101)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd102 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(102)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd103 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(103)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd104 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(104)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd105 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(105)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd106 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(106)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd107 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(107)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd108 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(108)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd109 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(109)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd110 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(110)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd111 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(111)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd112 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(112)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd113 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(113)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd114 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(114)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd115 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(115)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd116 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(116)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd117 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(117)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd118 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(118)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd119 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(119)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd120 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(120)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd121 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(121)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd122 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(122)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd123 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(123)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd124 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(124)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd125 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(125)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd126 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(126)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd127 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(127)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd128 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(128)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd129 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(129)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd130 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(130)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd131 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(131)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd132 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(132)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd133 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(133)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd134 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(134)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd135 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(135)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd136 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(136)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd137 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(137)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd138 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(138)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd139 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(139)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd140 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(140)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd141 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(141)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd142 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(142)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd143 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(143)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd144 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(144)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd145 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(145)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd146 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(146)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd147 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(147)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd148 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(148)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd149 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(149)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd150 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(150)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd151 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(151)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd152 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(152)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd153 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(153)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd154 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(154)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd155 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(155)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd156 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(156)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd157 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(157)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd158 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(158)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd159 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(159)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd160 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(160)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd161 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(161)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd162 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(162)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd163 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(163)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd164 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(164)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd165 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(165)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd166 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(166)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd167 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(167)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd168 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(168)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd169 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(169)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd170 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(170)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd171 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(171)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd172 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(172)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd173 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(173)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd174 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(174)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd175 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(175)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd176 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(176)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd177 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(177)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd178 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(178)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd179 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(179)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd180 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(180)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd181 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(181)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd182 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(182)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd183 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(183)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd184 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(184)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd185 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(185)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd186 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(186)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd187 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(187)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd188 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(188)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd189 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(189)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd190 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(190)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd191 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(191)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd192 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(192)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd193 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(193)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd194 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(194)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd195 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(195)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd196 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(196)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd197 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(197)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd198 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(198)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd199 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(199)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd200 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(200)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd201 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(201)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd202 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(202)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd203 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(203)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd204 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(204)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd205 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(205)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd206 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(206)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd207 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(207)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd208 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(208)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd209 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(209)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd210 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(210)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd211 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(211)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd212 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(212)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd213 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(213)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd214 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(214)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd215 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(215)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd216 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(216)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd217 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(217)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd218 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(218)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd219 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(219)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd220 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(220)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd221 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(221)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd222 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(222)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd223 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(223)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd224 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(224)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd225 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(225)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd226 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(226)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd227 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(227)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd228 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(228)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd229 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(229)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd230 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(230)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd231 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(231)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd232 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(232)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd233 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(233)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd234 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(234)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd235 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(235)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd236 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(236)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd237 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(237)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd238 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(238)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd239 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(239)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd240 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(240)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd241 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(241)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd242 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(242)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd243 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(243)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd244 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(244)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd245 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(245)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd246 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(246)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd247 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(247)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd248 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(248)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd249 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(249)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd250 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(250)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd251 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(251)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd252 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(252)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd253 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(253)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd254 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(254)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd255 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(255)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd256 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(256)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd257 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(257)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd258 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(258)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd259 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(259)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd260 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(260)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd261 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(261)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd262 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(262)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd263 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(263)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd264 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(264)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd265 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(265)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd266 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(266)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd267 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(267)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd268 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(268)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd269 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(269)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd270 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(270)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd271 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(271)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd272 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(272)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd273 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(273)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd274 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(274)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd275 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(275)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd276 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(276)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd277 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(277)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd278 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(278)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd279 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(279)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd280 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(280)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd281 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(281)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd282 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(282)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd283 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(283)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd284 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(284)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd285 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(285)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd286 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(286)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd287 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(287)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd288 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(288)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd289 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(289)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd290 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(290)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd291 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(291)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd292 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(292)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd293 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(293)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd294 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(294)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd295 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(295)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd296 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(296)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd297 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(297)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd298 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(298)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd299 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(299)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd300 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(300)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd301 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(301)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd302 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(302)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd303 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(303)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd304 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(304)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd305 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(305)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd306 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(306)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd307 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(307)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd308 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(308)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd309 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(309)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd310 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(310)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd311 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(311)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd312 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(312)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd313 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(313)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd314 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(314)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd315 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(315)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd316 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(316)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd317 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(317)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd318 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(318)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd319 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(319)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd320 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(320)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd321 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(321)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd322 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(322)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd323 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(323)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd324 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(324)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd325 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(325)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd326 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(326)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd327 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(327)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd328 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(328)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd329 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(329)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd330 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(330)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd331 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(331)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd332 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(332)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd333 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(333)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd334 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(334)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd335 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(335)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd336 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(336)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd337 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(337)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd338 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(338)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd339 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(339)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd340 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(340)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd341 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(341)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd342 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(342)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd343 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(343)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd344 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(344)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd345 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(345)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd346 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(346)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd347 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(347)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd348 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(348)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd349 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(349)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd350 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(350)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd351 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(351)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd352 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(352)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd353 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(353)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd354 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(354)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd355 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(355)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd356 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(356)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd357 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(357)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd358 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(358)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd359 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(359)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd360 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(360)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd361 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(361)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd362 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(362)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd363 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(363)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd364 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(364)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd365 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(365)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd366 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(366)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd367 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(367)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd368 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(368)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd369 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(369)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd370 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(370)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd371 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(371)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd372 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(372)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd373 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(373)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd374 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(374)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd375 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(375)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd376 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(376)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd377 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(377)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd378 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(378)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd379 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(379)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd380 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(380)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd381 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(381)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd382 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(382)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd383 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(383)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd384 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(384)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd385 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(385)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd386 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(386)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd387 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(387)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd388 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(388)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd389 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(389)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd390 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(390)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd391 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(391)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd392 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(392)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd393 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(393)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd394 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(394)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd395 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(395)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd396 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(396)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd397 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(397)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd398 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(398)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd399 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(399)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd400 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(400)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd401 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(401)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd402 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(402)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd403 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(403)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd404 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(404)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd405 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(405)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd406 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(406)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd407 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(407)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd408 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(408)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd409 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(409)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd410 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(410)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd411 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(411)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd412 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(412)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd413 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(413)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd414 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(414)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd415 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(415)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd416 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(416)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd417 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(417)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd418 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(418)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd419 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(419)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd420 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(420)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd421 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(421)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd422 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(422)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd423 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(423)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd424 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(424)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd425 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(425)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd426 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(426)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd427 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(427)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd428 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(428)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd429 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(429)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd430 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(430)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd431 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(431)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd432 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(432)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd433 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(433)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd434 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(434)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd435 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(435)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd436 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(436)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd437 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(437)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd438 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(438)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd439 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(439)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd440 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(440)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd441 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(441)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd442 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(442)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd443 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(443)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd444 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(444)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd445 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(445)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd446 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(446)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd447 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(447)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd448 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(448)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd449 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(449)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd450 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(450)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd451 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(451)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd452 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(452)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd453 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(453)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd454 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(454)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd455 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(455)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd456 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(456)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd457 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(457)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd458 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(458)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd459 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(459)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd460 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(460)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd461 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(461)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd462 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(462)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd463 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(463)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd464 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(464)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd465 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(465)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd466 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(466)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd467 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(467)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd468 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(468)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd469 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(469)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd470 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(470)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd471 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(471)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd472 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(472)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd473 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(473)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd474 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(474)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd475 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(475)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd476 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(476)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd477 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(477)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd478 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(478)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd479 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(479)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd480 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(480)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd481 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(481)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd482 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(482)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd483 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(483)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd484 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(484)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd485 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(485)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd486 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(486)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd487 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(487)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd488 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(488)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd489 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(489)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd490 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(490)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd491 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(491)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd492 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(492)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd493 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(493)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd494 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(494)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd495 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(495)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd496 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(496)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd497 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(497)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd498 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(498)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd499 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(499)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd500 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(500)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd501 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(501)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd502 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(502)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd503 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(503)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd504 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(504)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd505 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(505)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd506 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(506)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd507 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(507)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd508 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(508)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd509 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(509)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd510 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(510)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd511 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(511)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd512 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(512)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd513 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(513)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd514 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(514)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd515 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(515)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd516 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(516)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd517 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(517)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd518 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(518)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd519 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(519)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd520 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(520)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd521 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(521)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd522 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(522)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd523 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(523)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd524 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(524)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd525 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(525)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd526 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(526)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd527 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(527)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd528 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(528)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd529 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(529)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd530 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(530)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd531 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(531)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd532 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(532)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd533 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(533)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd534 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(534)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd535 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(535)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd536 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(536)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd537 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(537)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd538 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(538)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd539 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(539)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd540 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(540)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd541 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(541)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd542 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(542)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd543 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(543)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd544 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(544)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd545 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(545)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd546 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(546)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd547 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(547)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd548 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(548)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd549 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(549)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd550 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(550)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd551 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(551)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd552 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(552)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd553 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(553)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd554 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(554)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd555 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(555)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd556 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(556)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd557 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(557)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd558 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(558)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd559 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(559)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd560 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(560)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd561 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(561)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd562 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(562)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd563 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(563)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd564 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(564)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd565 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(565)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd566 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(566)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd567 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(567)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd568 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(568)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd569 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(569)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd570 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(570)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd571 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(571)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd572 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(572)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd573 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(573)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd574 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(574)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd575 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(575)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd576 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(576)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd577 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(577)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd578 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(578)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd579 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(579)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd580 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(580)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd581 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(581)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd582 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(582)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd583 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(583)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd584 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(584)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd585 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(585)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd586 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(586)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd587 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(587)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd588 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(588)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd589 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(589)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd590 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(590)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd591 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(591)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd592 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(592)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd593 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(593)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd594 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(594)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd595 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(595)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd596 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(596)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd597 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(597)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd598 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(598)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd599 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(599)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd600 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(600)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd601 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(601)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd602 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(602)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd603 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(603)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd604 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(604)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd605 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(605)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd606 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(606)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd607 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(607)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd608 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(608)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd609 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(609)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd610 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(610)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd611 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(611)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd612 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(612)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd613 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(613)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd614 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(614)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd615 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(615)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd616 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(616)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd617 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(617)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd618 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(618)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd619 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(619)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd620 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(620)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd621 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(621)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd622 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(622)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd623 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(623)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd624 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(624)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd625 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(625)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd626 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(626)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd627 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(627)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd628 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(628)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd629 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(629)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd630 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(630)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd631 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(631)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd632 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(632)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd633 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(633)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd634 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(634)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd635 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(635)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd636 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(636)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd637 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(637)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd638 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(638)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd639 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(639)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd640 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(640)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd641 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(641)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd642 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(642)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd643 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(643)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd644 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(644)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd645 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(645)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd646 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(646)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd647 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(647)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd648 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(648)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd649 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(649)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd650 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(650)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd651 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(651)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd652 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(652)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd653 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(653)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd654 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(654)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd655 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(655)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd656 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(656)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd657 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(657)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd658 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(658)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd659 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(659)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd660 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(660)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd661 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(661)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd662 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(662)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd663 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(663)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd664 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(664)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd665 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(665)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd666 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(666)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd667 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(667)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd668 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(668)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd669 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(669)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd670 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(670)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd671 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(671)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd672 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(672)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd673 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(673)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd674 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(674)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd675 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(675)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd676 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(676)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd677 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(677)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd678 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(678)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd679 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(679)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd680 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(680)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd681 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(681)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd682 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(682)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd683 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(683)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd684 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(684)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd685 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(685)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd686 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(686)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd687 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(687)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd688 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(688)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd689 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(689)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd690 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(690)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd691 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(691)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd692 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(692)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd693 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(693)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd694 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(694)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd695 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(695)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd696 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(696)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd697 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(697)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd698 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(698)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd699 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(699)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd700 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(700)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd701 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(701)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd702 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(702)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd703 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(703)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd704 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(704)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd705 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(705)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd706 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(706)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd707 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(707)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd708 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(708)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd709 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(709)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd710 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(710)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd711 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(711)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd712 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(712)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd713 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(713)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd714 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(714)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd715 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(715)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd716 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(716)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd717 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(717)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd718 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(718)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd719 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(719)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd720 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(720)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd721 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(721)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd722 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(722)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd723 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(723)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd724 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(724)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd725 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(725)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd726 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(726)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd727 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(727)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd728 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(728)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd729 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(729)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd730 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(730)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd731 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(731)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd732 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(732)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd733 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(733)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd734 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(734)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd735 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(735)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd736 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(736)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd737 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(737)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd738 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(738)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd739 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(739)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd740 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(740)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd741 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(741)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd742 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(742)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd743 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(743)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd744 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(744)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd745 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(745)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd746 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(746)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd747 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(747)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd748 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(748)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd749 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(749)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd750 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(750)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd751 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(751)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd752 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(752)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd753 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(753)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd754 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(754)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd755 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(755)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd756 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(756)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd757 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(757)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd758 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(758)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd759 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(759)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd760 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(760)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd761 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(761)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd762 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(762)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd763 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(763)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd764 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(764)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd765 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(765)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd766 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(766)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd767 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(767)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd768 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(768)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd769 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(769)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd770 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(770)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd771 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(771)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd772 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(772)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd773 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(773)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd774 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(774)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd775 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(775)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd776 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(776)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd777 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(777)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd778 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(778)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd779 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(779)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd780 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(780)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd781 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(781)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd782 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(782)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd783 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(783)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd784 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(784)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd785 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(785)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd786 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(786)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd787 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(787)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd788 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(788)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd789 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(789)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd790 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(790)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd791 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(791)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd792 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(792)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd793 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(793)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd794 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(794)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd795 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(795)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd796 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(796)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd797 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(797)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd798 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(798)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd799 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(799)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd800 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(800)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd801 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(801)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd802 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(802)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd803 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(803)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd804 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(804)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd805 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(805)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd806 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(806)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd807 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(807)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd808 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(808)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd809 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(809)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd810 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(810)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd811 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(811)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd812 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(812)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd813 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(813)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd814 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(814)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd815 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(815)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd816 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(816)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd817 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(817)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd818 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(818)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd819 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(819)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd820 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(820)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd821 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(821)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd822 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(822)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd823 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(823)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd824 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(824)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd825 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(825)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd826 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(826)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd827 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(827)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd828 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(828)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd829 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(829)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd830 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(830)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd831 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(831)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd832 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(832)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd833 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(833)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd834 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(834)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd835 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(835)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd836 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(836)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd837 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(837)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd838 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(838)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd839 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(839)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd840 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(840)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd841 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(841)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd842 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(842)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd843 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(843)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd844 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(844)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd845 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(845)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd846 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(846)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd847 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(847)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd848 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(848)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd849 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(849)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd850 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(850)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd851 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(851)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd852 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(852)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd853 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(853)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd854 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(854)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd855 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(855)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd856 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(856)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd857 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(857)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd858 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(858)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd859 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(859)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd860 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(860)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd861 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(861)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd862 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(862)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd863 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(863)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd864 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(864)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd865 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(865)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd866 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(866)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd867 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(867)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd868 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(868)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd869 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(869)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd870 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(870)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd871 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(871)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd872 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(872)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd873 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(873)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd874 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(874)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd875 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(875)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd876 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(876)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd877 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(877)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd878 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(878)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd879 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(879)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd880 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(880)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd881 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(881)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd882 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(882)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd883 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(883)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd884 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(884)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd885 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(885)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd886 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(886)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd887 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(887)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd888 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(888)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd889 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(889)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd890 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(890)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd891 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(891)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd892 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(892)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd893 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(893)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd894 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(894)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd895 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(895)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd896 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(896)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd897 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(897)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd898 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(898)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd899 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(899)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd900 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(900)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd901 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(901)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd902 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(902)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd903 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(903)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd904 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(904)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd905 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(905)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd906 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(906)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd907 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(907)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd908 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(908)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd909 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(909)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd910 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(910)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd911 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(911)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd912 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(912)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd913 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(913)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd914 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(914)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd915 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(915)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd916 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(916)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd917 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(917)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd918 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(918)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd919 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(919)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd920 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(920)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd921 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(921)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd922 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(922)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd923 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(923)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd924 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(924)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd925 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(925)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd926 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(926)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd927 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(927)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd928 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(928)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd929 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(929)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd930 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(930)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd931 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(931)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd932 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(932)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd933 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(933)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd934 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(934)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd935 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(935)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd936 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(936)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd937 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(937)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd938 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(938)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd939 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(939)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd940 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(940)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd941 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(941)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd942 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(942)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd943 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(943)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd944 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(944)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd945 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(945)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd946 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(946)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd947 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(947)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd948 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(948)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd949 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(949)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd950 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(950)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd951 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(951)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd952 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(952)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd953 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(953)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd954 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(954)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd955 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(955)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd956 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(956)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd957 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(957)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd958 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(958)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd959 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(959)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd960 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(960)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd961 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(961)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd962 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(962)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd963 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(963)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd964 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(964)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd965 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(965)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd966 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(966)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd967 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(967)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd968 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(968)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd969 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(969)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd970 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(970)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd971 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(971)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd972 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(972)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd973 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(973)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd974 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(974)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd975 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(975)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd976 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(976)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd977 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(977)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd978 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(978)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd979 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(979)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd980 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(980)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd981 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(981)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd982 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(982)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd983 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(983)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd984 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(984)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd985 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(985)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd986 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(986)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd987 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(987)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd988 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(988)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd989 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(989)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd990 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(990)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd991 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(991)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd992 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(992)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd993 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(993)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd994 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(994)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd995 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(995)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd996 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(996)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd997 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(997)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd998 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(998)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd999 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(999)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1000 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1000)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1001 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1001)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1002 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1002)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1003 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1003)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1004 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1004)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1005 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1005)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1006 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1006)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1007 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1007)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1008 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1008)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1009 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1009)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1010 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1010)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1011 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1011)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1012 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1012)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1013 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1013)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1014 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1014)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1015 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1015)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1016 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1016)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1017 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1017)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1018 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1018)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1019 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1019)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1020 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1020)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1021 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1021)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1022 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1022)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1023 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1023)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1024 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1024)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1025 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1025)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1026 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1026)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1027 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1027)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1028 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1028)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1029 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1029)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1030 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1030)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1031 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1031)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1032 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1032)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1033 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1033)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1034 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1034)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1035 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1035)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1036 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1036)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1037 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1037)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1038 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1038)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1039 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1039)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1040 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1040)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1041 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1041)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1042 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1042)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1043 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1043)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1044 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1044)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1045 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1045)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1046 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1046)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1047 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1047)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1048 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1048, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1048)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1049 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1049, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1049)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1050 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1050, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1050)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1051 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1051, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1051)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1052 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1052, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1052)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1053 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1053, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1053)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1054 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1054, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1054)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1055 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1055, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1055)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1056 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1056, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1056)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1057 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1057, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1057)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1058 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1058, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1058)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1059 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1059, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1059)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1060 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1060, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1060)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1061 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1061, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1061)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1062 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1062, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1062)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1063 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1063, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1063)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1064 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1064, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1064)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1065 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1065, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1065)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1066 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1066, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1066)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1067 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1067, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1067)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1068 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1068, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1068)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1069 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1069, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1069)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1070 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1070, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1070)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1071 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1071, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1071)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1072 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1072, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1072)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1073 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1073, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1073)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1074 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1074, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1074)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1075 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1075, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1075)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1076 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1076, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1076)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1077 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1077, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1077)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1078 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1078, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1078)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1079 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1079, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1079)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1080 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1080, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1080)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1081 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1081, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1081)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1082 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1082, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1082)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1083 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1083, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1083)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1084 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1084, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1084)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1085 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1085, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1085)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1086 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1086, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1086)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1087 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1087, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1087)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1088 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1088, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1088)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1089 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1089, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1089)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1090 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1090, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1090)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1091 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1091, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1091)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1092 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1092, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1092)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1093 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1093, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1093)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1094 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1094, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1094)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1095 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1095, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1095)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1096 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1096, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1096)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1097 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1097, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1097)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1098 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1098, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1098)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1099 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1099, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1099)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1100 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1100, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1100)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1101 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1101, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1101)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1102 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1102, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1102)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1103 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1103, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1103)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1104 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1104, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1104)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1105 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1105, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1105)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1106 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1106, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1106)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1107 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1107, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1107)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1108 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1108, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1108)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1109 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1109, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1109)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1110 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1110, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1110)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1111 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1111, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1111)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1112 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1112, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1112)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1113 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1113, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1113)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1114 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1114, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1114)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1115 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1115, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1115)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1116 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1116, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1116)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1117 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1117, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1117)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1118 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1118, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1118)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1119 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1119, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1119)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1120 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1120, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1120)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1121 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1121, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1121)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1122 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1122, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1122)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1123 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1123, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1123)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1124 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1124, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1124)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1125 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1125, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1125)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1126 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1126, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1126)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1127 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1127, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1127)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1128 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1128, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1128)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1129 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1129, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1129)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1130 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1130, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1130)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1131 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1131, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1131)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1132 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1132, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1132)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1133 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1133, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1133)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1134 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1134, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1134)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1135 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1135, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1135)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1136 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1136, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1136)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1137 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1137, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1137)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1138 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1138, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1138)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1139 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1139, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1139)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1140 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1140, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1140)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1141 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1141, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1141)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1142 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1142, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1142)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1143 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1143, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1143)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1144 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1144, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1144)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1145 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1145, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1145)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1146 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1146, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1146)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1147 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1147, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1147)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1148 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1148, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1148)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1149 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1149, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1149)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1150 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1150, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1150)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1151 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1151, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1151)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1152 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1152, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1152)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1153 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1153, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1153)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1154 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1154, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1154)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1155 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1155, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1155)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1156 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1156, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1156)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1157 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1157, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1157)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1158 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1158, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1158)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1159 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1159, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1159)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1160 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1160, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1160)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1161 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1161, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1161)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1162 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1162, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1162)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1163 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1163, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1163)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1164 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1164, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1164)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1165 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1165, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1165)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1166 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1166, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1166)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1167 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1167, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1167)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1168 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1168, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1168)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1169 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1169, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1169)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1170 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1170, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1170)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1171 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1171, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1171)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1172 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1172, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1172)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1173 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1173, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1173)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1174 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1174, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1174)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1175 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1175, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1175)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1176 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1176, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1176)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1177 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1177, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1177)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1178 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1178, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1178)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1179 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1179, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1179)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1180 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1180, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1180)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1181 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1181, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1181)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1182 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1182, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1182)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1183 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1183, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1183)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1184 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1184, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1184)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1185 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1185, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1185)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1186 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1186, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1186)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1187 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1187, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1187)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1188 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1188, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1188)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1189 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1189, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1189)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1190 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1190, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1190)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1191 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1191, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1191)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1192 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1192, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1192)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1193 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1193, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1193)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1194 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1194, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1194)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1195 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1195, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1195)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1196 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1196, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1196)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1197 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1197, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1197)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1198 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1198, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1198)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1199 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1199, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1199)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1200 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1200, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1200)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1201 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1201, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1201)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1202 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1202, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1202)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1203 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1203, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1203)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1204 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1204, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1204)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1205 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1205, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1205)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1206 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1206, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1206)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1207 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1207, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1207)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1208 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1208, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1208)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1209 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1209, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1209)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1210 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1210, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1210)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1211 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1211, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1211)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1212 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1212, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1212)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1213 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1213, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1213)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1214 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1214, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1214)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1215 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1215, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1215)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1216 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1216, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1216)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1217 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1217, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1217)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1218 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1218, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1218)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1219 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1219, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1219)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1220 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1220, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1220)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1221 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1221, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1221)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1222 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1222, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1222)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1223 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1223, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1223)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1224 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1224, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1224)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1225 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1225, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1225)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1226 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1226, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1226)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1227 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1227, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1227)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1228 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1228, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1228)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1229 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1229, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1229)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1230 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1230, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1230)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1231 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1231, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1231)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1232 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1232, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1232)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1233 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1233, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1233)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1234 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1234, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1234)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1235 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1235, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1235)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1236 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1236, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1236)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1237 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1237, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1237)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1238 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1238, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1238)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1239 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1239, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1239)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1240 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1240, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1240)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1241 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1241, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1241)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1242 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1242, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1242)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1243 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1243, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1243)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1244 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1244, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1244)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1245 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1245, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1245)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1246 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1246, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1246)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1247 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1247, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1247)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1248 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1248, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1248)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1249 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1249, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1249)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1250 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1250, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1250)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1251 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1251, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1251)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1252 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1252, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1252)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1253 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1253, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1253)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1254 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1254, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1254)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1255 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1255, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1255)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1256 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1256, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1256)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1257 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1257, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1257)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1258 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1258, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1258)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1259 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1259, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1259)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1260 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1260, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1260)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1261 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1261, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1261)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1262 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1262, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1262)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1263 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1263, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1263)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1264 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1264, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1264)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1265 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1265, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1265)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1266 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1266, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1266)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1267 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1267, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1267)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1268 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1268, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1268)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1269 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1269, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1269)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1270 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1270, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1270)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1271 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1271, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1271)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1272 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1272, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1272)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1273 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1273, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1273)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1274 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1274, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1274)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1275 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1275, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1275)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1276 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1276, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1276)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1277 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1277, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1277)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1278 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1278, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1278)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1279 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1279, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1279)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1280 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1280, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1280)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1281 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1281, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1281)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1282 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1282, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1282)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1283 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1283, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1283)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1284 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1284, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1284)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1285 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1285, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1285)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1286 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1286, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1286)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1287 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1287, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1287)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1288 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1288, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1288)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1289 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1289, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1289)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1290 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1290, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1290)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1291 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1291, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1291)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1292 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1292, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1292)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1293 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1293, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1293)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1294 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1294, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1294)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1295 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1295, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1295)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1296 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1296, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1296)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1297 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1297, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1297)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1298 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1298, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1298)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1299 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1299, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1299)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1300 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1300, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1300)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1301 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1301, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1301)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1302 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1302, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1302)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1303 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1303, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1303)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1304 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1304, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1304)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1305 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1305, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1305)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1306 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1306, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1306)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1307 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1307, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1307)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1308 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1308, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1308)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1309 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1309, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1309)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1310 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1310, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1310)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1311 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1311, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1311)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1312 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1312, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1312)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1313 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1313, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1313)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1314 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1314, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1314)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1315 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1315, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1315)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1316 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1316, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1316)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1317 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1317, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1317)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1318 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1318, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1318)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1319 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1319, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1319)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1320 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1320, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1320)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1321 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1321, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1321)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1322 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1322, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1322)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1323 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1323, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1323)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1324 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1324, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1324)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1325 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1325, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1325)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1326 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1326, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1326)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1327 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1327, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1327)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1328 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1328, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1328)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1329 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1329, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1329)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1330 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1330, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1330)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1331 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1331, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1331)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1332 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1332, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1332)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1333 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1333, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1333)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1334 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1334, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1334)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1335 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1335, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1335)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1336 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1336, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1336)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1337 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1337, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1337)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1338 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1338, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1338)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1339 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1339, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1339)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1340 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1340, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1340)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1341 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1341, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1341)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1342 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1342, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1342)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1343 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1343, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1343)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1344 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1344, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1344)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1345 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1345, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1345)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1346 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1346, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1346)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1347 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1347, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1347)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1348 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1348, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1348)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1349 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1349, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1349)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1350 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1350, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1350)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1351 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1351, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1351)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1352 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1352, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1352)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1353 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1353, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1353)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1354 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1354, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1354)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1355 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1355, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1355)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1356 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1356, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1356)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1357 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1357, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1357)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1358 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1358, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1358)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1359 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1359, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1359)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1360 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1360, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1360)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1361 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1361, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1361)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1362 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1362, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1362)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1363 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1363, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1363)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1364 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1364, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1364)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1365 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1365, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1365)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1366 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1366, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1366)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1367 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1367, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1367)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1368 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1368, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1368)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1369 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1369, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1369)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1370 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1370, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1370)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1371 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1371, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1371)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1372 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1372, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1372)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1373 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1373, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1373)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1374 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1374, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1374)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1375 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1375, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1375)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1376 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1376, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1376)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1377 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1377, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1377)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1378 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1378, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1378)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1379 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1379, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1379)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1380 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1380, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1380)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1381 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1381, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1381)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1382 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1382, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1382)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1383 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1383, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1383)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1384 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1384, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1384)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1385 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1385, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1385)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1386 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1386, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1386)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1387 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1387, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1387)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1388 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1388, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1388)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1389 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1389, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1389)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1390 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1390, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1390)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1391 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1391, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1391)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1392 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1392, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1392)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1393 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1393, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1393)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1394 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1394, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1394)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1395 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1395, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1395)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1396 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1396, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1396)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1397 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1397, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1397)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1398 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1398, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1398)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1399 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1399, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1399)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1400 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1400, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1400)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1401 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1401, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1401)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1402 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1402, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1402)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1403 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1403, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1403)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1404 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1404, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1404)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1405 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1405, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1405)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1406 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1406, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1406)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1407 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1407, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1407)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1408 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1408, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1408)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1409 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1409, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1409)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1410 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1410, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1410)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1411 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1411, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1411)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1412 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1412, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1412)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1413 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1413, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1413)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1414 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1414, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1414)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1415 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1415, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1415)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1416 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1416, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1416)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1417 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1417, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1417)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1418 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1418, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1418)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1419 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1419, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1419)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1420 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1420, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1420)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1421 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1421, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1421)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1422 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1422, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1422)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1423 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1423, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1423)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1424 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1424, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1424)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1425 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1425, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1425)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1426 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1426, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1426)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1427 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1427, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1427)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1428 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1428, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1428)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1429 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1429, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1429)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1430 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1430, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1430)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1431 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1431, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1431)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1432 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1432, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1432)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1433 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1433, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1433)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1434 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1434, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1434)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1435 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1435, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1435)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1436 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1436, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1436)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1437 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1437, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1437)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1438 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1438, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1438)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1439 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1439, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1439)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1440 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1440, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1440)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1441 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1441, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1441)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1442 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1442, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1442)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1443 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1443, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1443)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1444 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1444, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1444)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1445 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1445, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1445)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1446 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1446, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1446)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1447 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1447, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1447)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1448 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1448, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1448)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1449 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1449, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1449)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1450 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1450, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1450)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1451 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1451, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1451)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1452 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1452, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1452)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1453 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1453, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1453)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1454 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1454, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1454)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1455 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1455, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1455)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1456 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1456, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1456)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1457 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1457, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1457)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1458 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1458, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1458)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1459 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1459, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1459)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1460 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1460, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1460)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1461 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1461, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1461)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1462 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1462, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1462)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1463 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1463, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1463)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1464 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1464, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1464)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1465 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1465, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1465)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1466 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1466, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1466)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1467 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1467, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1467)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1468 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1468, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1468)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1469 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1469, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1469)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1470 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1470, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1470)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1471 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1471, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1471)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1472 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1472, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1472)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1473 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1473, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1473)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1474 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1474, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1474)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1475 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1475, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1475)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1476 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1476, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1476)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1477 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1477, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1477)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1478 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1478, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1478)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1479 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1479, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1479)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1480 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1480, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1480)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1481 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1481, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1481)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1482 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1482, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1482)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1483 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1483, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1483)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1484 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1484, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1484)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1485 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1485, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1485)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1486 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1486, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1486)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1487 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1487, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1487)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1488 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1488, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1488)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1489 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1489, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1489)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1490 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1490, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1490)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1491 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1491, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1491)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1492 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1492, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1492)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1493 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1493, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1493)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1494 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1494, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1494)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1495 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1495, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1495)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1496 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1496, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1496)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1497 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1497, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1497)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1498 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1498, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1498)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1499 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1499, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1499)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1500 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1500, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1500)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1501 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1501, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1501)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1502 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1502, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1502)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1503 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1503, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1503)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1504 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1504, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1504)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1505 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1505, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1505)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1506 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1506, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1506)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1507 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1507, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1507)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1508 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1508, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1508)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1509 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1509, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1509)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1510 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1510, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1510)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1511 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1511, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1511)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1512 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1512, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1512)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1513 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1513, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1513)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1514 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1514, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1514)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1515 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1515, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1515)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1516 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1516, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1516)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1517 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1517, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1517)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1518 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1518, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1518)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1519 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1519, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1519)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1520 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1520, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1520)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1521 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1521, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1521)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1522 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1522, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1522)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1523 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1523, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1523)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1524 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1524, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1524)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1525 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1525, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1525)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1526 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1526, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1526)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1527 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1527, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1527)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1528 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1528, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1528)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1529 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1529, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1529)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1530 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1530, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1530)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1531 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1531, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1531)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1532 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1532, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1532)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1533 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1533, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1533)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1534 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1534, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1534)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1535 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1535, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1535)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1536 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1536, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1536)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1537 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1537, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1537)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1538 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1538, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1538)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1539 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1539, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1539)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1540 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1540, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1540)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1541 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1541, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1541)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1542 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1542, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1542)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1543 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1543, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1543)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1544 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1544, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1544)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1545 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1545, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1545)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1546 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1546, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1546)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1547 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1547, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1547)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1548 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1548, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1548)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1549 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1549, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1549)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1550 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1550, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1550)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1551 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1551, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1551)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1552 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1552, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1552)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1553 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1553, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1553)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1554 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1554, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1554)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1555 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1555, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1555)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1556 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1556, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1556)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1557 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1557, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1557)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1558 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1558, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1558)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1559 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1559, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1559)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1560 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1560, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1560)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1561 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1561, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1561)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1562 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1562, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1562)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1563 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1563, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1563)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1564 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1564, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1564)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1565 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1565, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1565)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1566 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1566, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1566)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1567 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1567, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1567)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1568 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1568, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1568)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1569 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1569, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1569)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1570 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1570, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1570)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1571 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1571, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1571)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1572 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1572, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1572)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1573 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1573, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1573)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1574 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1574, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1574)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1575 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1575, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1575)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1576 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1576, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1576)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1577 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1577, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1577)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1578 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1578, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1578)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1579 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1579, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1579)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1580 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1580, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1580)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1581 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1581, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1581)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1582 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1582, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1582)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1583 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1583, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1583)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1584 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1584, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1584)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1585 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1585, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1585)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1586 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1586, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1586)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1587 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1587, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1587)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1588 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1588, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1588)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1589 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1589, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1589)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1590 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1590, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1590)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1591 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1591, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1591)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1592 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1592, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1592)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1593 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1593, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1593)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1594 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1594, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1594)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1595 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1595, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1595)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1596 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1596, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1596)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1597 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1597, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1597)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1598 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1598, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1598)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1599 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1599, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1599)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1600 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1600, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1600)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1601 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1601, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1601)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1602 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1602, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1602)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1603 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1603, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1603)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1604 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1604, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1604)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1605 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1605, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1605)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1606 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1606, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1606)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1607 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1607, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1607)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1608 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1608, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1608)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1609 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1609, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1609)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1610 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1610, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1610)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1611 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1611, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1611)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1612 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1612, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1612)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1613 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1613, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1613)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1614 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1614, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1614)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1615 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1615, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1615)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1616 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1616, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1616)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1617 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1617, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1617)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1618 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1618, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1618)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1619 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1619, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1619)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1620 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1620, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1620)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1621 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1621, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1621)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1622 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1622, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1622)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1623 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1623, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1623)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1624 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1624, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1624)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1625 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1625, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1625)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1626 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1626, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1626)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1627 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1627, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1627)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1628 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1628, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1628)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1629 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1629, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1629)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1630 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1630, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1630)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1631 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1631, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1631)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1632 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1632, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1632)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1633 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1633, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1633)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1634 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1634, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1634)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1635 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1635, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1635)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1636 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1636, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1636)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1637 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1637, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1637)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1638 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1638, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1638)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1639 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1639, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1639)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1640 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1640, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1640)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1641 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1641, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1641)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1642 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1642, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1642)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1643 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1643, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1643)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1644 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1644, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1644)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1645 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1645, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1645)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1646 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1646, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1646)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1647 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1647, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1647)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1648 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1648, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1648)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1649 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1649, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1649)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1650 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1650, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1650)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1651 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1651, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1651)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1652 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1652, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1652)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1653 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1653, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1653)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1654 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1654, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1654)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1655 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1655, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1655)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1656 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1656, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1656)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1657 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1657, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1657)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1658 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1658, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1658)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1659 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1659, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1659)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1660 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1660, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1660)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1661 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1661, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1661)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1662 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1662, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1662)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1663 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1663, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1663)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1664 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1664, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1664)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1665 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1665, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1665)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1666 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1666, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1666)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1667 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1667, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1667)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1668 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1668, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1668)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1669 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1669, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1669)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1670 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1670, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1670)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1671 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1671, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1671)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1672 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1672, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1672)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1673 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1673, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1673)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1674 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1674, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1674)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1675 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1675, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1675)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1676 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1676, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1676)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1677 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1677, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1677)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1678 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1678, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1678)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1679 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1679, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1679)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1680 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1680, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1680)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1681 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1681, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1681)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1682 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1682, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1682)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1683 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1683, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1683)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1684 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1684, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1684)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1685 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1685, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1685)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1686 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1686, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1686)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1687 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1687, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1687)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1688 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1688, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1688)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1689 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1689, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1689)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1690 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1690, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1690)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1691 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1691, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1691)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1692 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1692, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1692)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1693 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1693, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1693)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1694 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1694, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1694)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1695 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1695, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1695)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1696 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1696, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1696)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1697 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1697, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1697)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1698 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1698, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1698)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1699 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1699, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1699)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1700 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1700, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1700)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1701 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1701, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1701)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1702 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1702, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1702)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1703 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1703, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1703)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1704 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1704, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1704)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1705 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1705, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1705)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1706 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1706, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1706)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1707 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1707, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1707)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1708 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1708, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1708)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1709 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1709, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1709)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1710 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1710, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1710)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1711 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1711, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1711)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1712 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1712, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1712)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1713 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1713, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1713)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1714 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1714, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1714)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1715 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1715, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1715)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1716 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1716, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1716)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1717 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1717, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1717)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1718 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1718, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1718)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1719 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1719, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1719)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1720 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1720, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1720)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1721 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1721, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1721)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1722 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1722, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1722)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1723 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1723, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1723)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1724 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1724, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1724)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1725 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1725, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1725)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1726 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1726, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1726)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1727 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1727, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1727)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1728 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1728, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1728)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1729 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1729, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1729)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1730 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1730, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1730)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1731 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1731, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1731)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1732 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1732, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1732)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1733 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1733, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1733)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1734 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1734, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1734)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1735 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1735, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1735)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1736 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1736, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1736)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1737 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1737, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1737)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1738 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1738, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1738)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1739 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1739, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1739)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1740 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1740, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1740)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1741 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1741, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1741)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1742 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1742, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1742)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1743 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1743, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1743)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1744 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1744, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1744)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1745 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1745, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1745)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1746 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1746, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1746)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1747 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1747, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1747)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1748 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1748, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1748)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1749 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1749, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1749)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1750 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1750, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1750)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1751 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1751, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1751)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1752 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1752, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1752)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1753 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1753, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1753)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1754 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1754, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1754)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1755 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1755, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1755)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1756 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1756, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1756)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1757 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1757, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1757)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1758 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1758, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1758)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1759 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1759, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1759)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1760 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1760, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1760)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1761 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1761, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1761)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1762 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1762, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1762)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1763 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1763, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1763)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1764 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1764, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1764)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1765 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1765, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1765)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1766 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1766, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1766)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1767 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1767, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1767)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1768 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1768, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1768)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1769 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1769, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1769)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1770 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1770, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1770)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1771 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1771, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1771)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1772 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1772, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1772)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1773 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1773, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1773)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1774 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1774, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1774)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1775 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1775, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1775)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1776 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1776, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1776)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1777 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1777, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1777)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1778 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1778, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1778)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1779 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1779, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1779)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1780 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1780, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1780)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1781 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1781, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1781)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1782 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1782, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1782)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1783 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1783, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1783)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1784 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1784, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1784)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1785 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1785, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1785)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1786 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1786, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1786)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1787 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1787, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1787)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1788 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1788, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1788)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1789 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1789, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1789)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1790 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1790, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1790)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1791 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1791, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1791)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1792 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1792, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1792)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1793 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1793, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1793)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1794 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1794, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1794)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1795 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1795, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1795)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1796 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1796, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1796)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1797 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1797, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1797)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1798 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1798, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1798)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1799 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1799, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1799)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1800 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1800, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1800)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1801 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1801, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1801)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1802 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1802, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1802)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1803 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1803, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1803)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1804 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1804, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1804)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1805 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1805, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1805)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1806 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1806, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1806)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1807 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1807, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1807)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1808 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1808, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1808)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1809 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1809, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1809)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1810 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1810, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1810)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1811 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1811, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1811)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1812 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1812, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1812)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1813 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1813, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1813)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1814 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1814, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1814)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1815 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1815, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1815)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1816 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1816, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1816)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1817 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1817, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1817)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1818 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1818, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1818)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1819 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1819, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1819)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1820 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1820, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1820)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1821 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1821, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1821)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1822 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1822, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1822)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1823 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1823, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1823)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1824 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1824, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1824)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1825 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1825, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1825)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1826 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1826, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1826)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1827 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1827, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1827)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1828 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1828, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1828)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1829 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1829, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1829)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1830 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1830, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1830)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1831 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1831, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1831)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1832 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1832, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1832)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1833 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1833, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1833)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1834 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1834, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1834)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1835 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1835, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1835)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1836 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1836, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1836)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1837 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1837, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1837)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1838 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1838, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1838)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1839 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1839, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1839)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1840 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1840, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1840)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1841 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1841, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1841)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1842 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1842, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1842)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1843 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1843, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1843)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1844 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1844, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1844)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1845 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1845, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1845)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1846 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1846, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1846)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1847 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1847, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1847)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1848 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1848, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1848)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1849 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1849, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1849)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1850 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1850, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1850)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1851 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1851, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1851)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1852 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1852, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1852)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1853 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1853, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1853)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1854 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1854, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1854)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1855 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1855, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1855)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1856 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1856, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1856)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1857 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1857, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1857)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1858 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1858, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1858)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1859 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1859, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1859)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1860 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1860, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1860)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1861 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1861, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1861)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1862 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1862, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1862)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1863 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1863, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1863)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1864 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1864, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1864)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1865 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1865, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1865)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1866 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1866, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1866)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1867 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1867, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1867)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1868 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1868, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1868)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1869 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1869, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1869)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1870 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1870, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1870)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1871 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1871, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1871)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1872 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1872, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1872)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1873 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1873, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1873)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1874 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1874, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1874)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1875 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1875, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1875)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1876 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1876, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1876)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1877 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1877, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1877)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1878 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1878, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1878)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1879 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1879, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1879)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1880 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1880, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1880)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1881 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1881, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1881)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1882 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1882, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1882)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1883 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1883, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1883)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1884 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1884, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1884)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1885 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1885, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1885)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1886 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1886, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1886)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1887 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1887, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1887)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1888 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1888, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1888)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1889 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1889, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1889)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1890 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1890, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1890)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1891 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1891, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1891)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1892 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1892, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1892)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1893 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1893, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1893)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1894 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1894, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1894)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1895 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1895, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1895)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1896 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1896, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1896)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1897 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1897, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1897)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1898 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1898, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1898)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1899 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1899, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1899)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1900 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1900, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1900)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1901 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1901, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1901)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1902 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1902, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1902)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1903 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1903, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1903)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1904 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1904, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1904)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1905 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1905, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1905)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1906 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1906, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1906)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1907 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1907, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1907)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1908 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1908, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1908)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1909 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1909, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1909)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1910 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1910, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1910)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1911 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1911, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1911)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1912 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1912, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1912)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1913 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1913, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1913)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1914 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1914, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1914)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1915 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1915, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1915)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1916 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1916, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1916)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1917 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1917, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1917)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1918 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1918, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1918)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1919 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1919, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1919)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1920 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1920, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1920)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1921 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1921, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1921)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1922 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1922, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1922)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1923 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1923, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1923)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1924 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1924, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1924)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1925 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1925, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1925)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1926 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1926, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1926)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1927 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1927, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1927)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1928 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1928, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1928)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1929 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1929, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1929)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1930 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1930, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1930)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1931 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1931, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1931)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1932 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1932, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1932)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1933 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1933, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1933)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1934 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1934, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1934)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1935 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1935, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1935)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1936 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1936, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1936)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1937 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1937, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1937)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1938 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1938, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1938)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1939 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1939, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1939)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1940 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1940, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1940)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1941 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1941, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1941)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1942 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1942, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1942)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1943 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1943, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1943)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1944 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1944, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1944)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1945 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1945, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1945)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1946 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1946, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1946)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1947 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1947, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1947)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1948 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1948, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1948)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1949 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1949, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1949)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1950 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1950, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1950)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1951 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1951, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1951)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1952 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1952, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1952)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1953 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1953, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1953)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1954 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1954, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1954)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1955 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1955, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1955)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1956 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1956, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1956)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1957 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1957, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1957)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1958 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1958, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1958)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1959 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1959, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1959)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1960 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1960, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1960)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1961 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1961, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1961)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1962 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1962, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1962)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1963 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1963, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1963)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1964 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1964, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1964)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1965 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1965, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1965)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1966 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1966, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1966)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1967 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1967, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1967)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1968 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1968, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1968)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1969 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1969, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1969)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1970 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1970, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1970)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1971 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1971, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1971)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1972 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1972, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1972)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1973 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1973, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1973)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1974 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1974, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1974)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1975 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1975, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1975)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1976 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1976, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1976)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1977 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1977, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1977)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1978 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1978, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1978)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1979 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1979, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1979)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1980 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1980, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1980)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1981 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1981, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1981)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1982 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1982, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1982)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1983 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1983, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1983)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1984 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1984, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1984)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1985 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1985, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1985)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1986 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1986, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1986)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1987 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1987, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1987)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1988 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1988, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1988)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1989 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1989, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1989)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1990 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1990, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1990)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1991 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1991, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1991)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1992 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1992, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1992)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1993 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1993, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1993)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1994 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1994, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1994)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1995 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1995, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1995)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1996 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1996, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1996)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1997 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1997, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1997)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1998 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1998, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1998)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd1999 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D1999, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(1999)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2000 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2000, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2000)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2001 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2001, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2001)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2002 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2002, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2002)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2003 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2003, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2003)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2004 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2004, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2004)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2005 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2005, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2005)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2006 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2006, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2006)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2007 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2007, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2007)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2008 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2008, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2008)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2009 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2009, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2009)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2010 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2010, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2010)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2011 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2011, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2011)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2012 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2012, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2012)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2013 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2013, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2013)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2014 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2014, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2014)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2015 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2015, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2015)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2016 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2016, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2016)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2017 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2017, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2017)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2018 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2018, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2018)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2019 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2019, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2019)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2020 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2020, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2020)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2021 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2021, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2021)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2022 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2022, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2022)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2023 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2023, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2023)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2024 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2024, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2024)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2025 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2025, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2025)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2026 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2026, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2026)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2027 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2027, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2027)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2028 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2028, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2028)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2029 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2029, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2029)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2030 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2030, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2030)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2031 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2031, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2031)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2032 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2032, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2032)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2033 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2033, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2033)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2034 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2034, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2034)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2035 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2035, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2035)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2036 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2036, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2036)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2037 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2037, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2037)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2038 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2038, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2038)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2039 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2039, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2039)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2040 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2040, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2040)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2041 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2041, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2041)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2042 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2042, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2042)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2043 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2043, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2043)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2044 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2044, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2044)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2045 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2045, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2045)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2046 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2046, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2046)
             
	end
         else if(local_pf_num == 'h0 && local_vf_num == 'd2047 && local_vf_active == 'h1) begin
          `uvm_do_on_with(master_seq, p_sequencer.master_sequencer_D2047, { tlp_length  == local_tlp_length  ;
                                                                         pf_num      == local_pf_num      ;
                                                                         vf_num      == local_vf_num      ;
                                                                         vf_active   == local_vf_active   ;
                                                                         payload     == local_payload     ;
                                                                         direction   == 1'b1              ;

                                                                        })

        `reset_in_middle(2047)
             
	end

