// Copyright (C) 2023 Intel Corporation
// SPDX-License-Identifier: MIT

/**
 * Abstract:
 * This file creates a basetest, which serves as the base class for the rest
 * of the tests in this environment.  This test sets up the default behavior
 * for the rest of the tests in this environment.
 *
 * In the build_phase phase of the test we will set the necessary test related 
 * information:
 *  - Create the pf_vf_mux_basic_env instance (named env)
 *  - Configure the pf_vf_mux_simple_reset_sequence as the default sequence
 *    for the reset phase of the TB ENV virtual sequencer
 */
`ifndef GUARD_PF_VF_MUX_BASE_TEST_SV
`define GUARD_PF_VF_MUX_BASE_TEST_SV

`include "pf_vf_mux_basic_env.sv"
`include "pf_vf_mux_simple_reset_sequence.sv"


class pf_vf_mux_base_test extends uvm_test;

  /** UVM Component Utility macro */
  `uvm_component_utils(pf_vf_mux_base_test)

  /** Instance of the environment */
  pf_vf_mux_basic_env env;
  int packet_count;

  //For stress_test
  int port_count[2048];

  /** Class Constructor */
  function new(string name = "pf_vf_mux_base_test", uvm_component parent=null);
    super.new(name,parent);
  endfunction: new

  /**
   * Build Phase
   * - Create the TB ENV
   * - Set the default sequences
   */

  virtual function void build_phase(uvm_phase phase);
    `uvm_info("build_phase", "Entered...", UVM_LOW)
    super.build_phase(phase);

    /** Create the environment */
    env = pf_vf_mux_basic_env::type_id::create("env", this);

    uvm_config_db#(uvm_object_wrapper)::set(this, "env.sequencer.reset_phase", "default_sequence", pf_vf_mux_simple_reset_sequence::type_id::get());

    `uvm_info("build_phase", "Exiting...", UVM_LOW)
  endfunction: build_phase


   function void end_of_elaboration_phase(uvm_phase phase);
    `SVT_XVM(root) root = `SVT_XVM(root)::get();
    uvm_object_wrapper _get_slave_resp_seq_item;
    `uvm_info("end_of_elaboration_phase", "Entered...", UVM_LOW)
   `uvm_info("BASE_TEST", "DISABLE_VIP_ERR ...",UVM_LOW)
    env.pf_vf_mux_system_env_H.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_H.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
    `ifdef TB_CONFIG_4
      env.pf_vf_mux_system_env_D.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      
      env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      
      env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif
    `ifdef TB_CONFIG_2
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif
    `ifdef TB_CONFIG_3
      env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif  

    env.pf_vf_mux_system_env_H.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_H.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[1].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[2].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[3].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[4].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[5].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[6].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[7].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[8].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[9].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[10].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[11].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[12].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[13].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[14].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[15].monitor.checks.signal_valid_tvalid_check);
    `ifdef TB_CONFIG_4
   env.pf_vf_mux_system_env_D.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[16].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[17].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[18].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[19].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[20].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[21].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[22].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[23].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[24].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[25].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[26].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[27].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[28].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[29].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[30].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[31].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[32].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[33].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[34].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[35].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[36].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[37].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[38].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[39].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[40].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[41].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[42].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[43].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[44].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[45].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[46].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[47].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[48].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[49].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[50].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[51].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[52].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[53].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[54].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[55].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[56].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[57].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[58].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[59].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[60].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[61].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[62].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[63].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[64].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[65].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[66].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[67].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[68].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[69].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[70].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[71].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[72].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[73].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[74].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[75].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[76].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[77].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[78].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[79].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[80].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[81].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[82].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[83].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[84].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[85].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[86].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[87].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[88].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[89].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[90].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[91].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[92].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[93].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[94].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[95].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[96].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[97].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[98].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[99].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[100].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[101].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[102].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[103].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[104].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[105].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[106].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[107].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[108].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[109].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[110].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[111].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[112].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[113].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[114].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[115].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[116].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[117].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[118].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[119].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[120].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[121].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[122].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[123].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[124].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[125].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[126].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[127].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[128].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[129].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[130].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[131].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[132].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[133].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[134].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[135].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[136].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[137].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[138].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[139].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[140].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[141].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[142].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[143].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[144].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[145].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[146].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[147].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[148].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[149].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[150].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[151].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[152].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[153].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[154].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[155].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[156].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[157].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[158].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[159].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[160].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[161].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[162].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[163].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[164].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[165].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[166].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[167].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[168].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[169].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[170].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[171].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[172].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[173].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[174].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[175].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[176].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[177].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[178].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[179].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[180].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[181].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[182].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[183].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[184].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[185].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[186].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[187].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[188].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[189].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[190].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[191].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[192].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[193].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[194].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[195].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[196].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[197].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[198].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[199].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[200].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[201].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[202].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[203].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[204].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[205].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[206].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[207].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[208].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[209].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[210].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[211].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[212].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[213].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[214].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[215].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[216].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[217].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[218].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[219].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[220].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[221].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[222].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[223].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[224].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[225].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[226].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[227].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[228].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[229].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[230].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[231].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[232].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[233].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[234].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[235].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[236].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[237].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[238].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[239].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[240].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[241].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[242].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[243].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[244].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[245].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[246].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[247].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[248].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[249].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[250].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[251].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[252].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[253].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[254].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[255].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[256].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[257].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[258].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[259].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[260].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[261].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[262].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[263].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[264].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[265].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[266].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[267].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[268].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[269].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[270].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[271].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[272].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[273].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[274].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[275].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[276].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[277].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[278].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[279].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[280].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[281].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[282].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[283].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[284].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[285].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[286].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[287].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[288].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[289].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[290].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[291].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[292].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[293].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[294].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[295].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[296].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[297].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[298].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[299].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[300].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[301].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[302].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[303].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[304].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[305].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[306].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[307].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[308].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[309].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[310].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[311].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[312].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[313].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[314].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[315].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[316].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[317].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[318].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[319].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[320].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[321].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[322].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[323].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[324].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[325].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[326].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[327].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[328].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[329].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[330].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[331].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[332].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[333].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[334].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[335].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[336].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[337].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[338].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[339].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[340].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[341].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[342].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[343].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[344].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[345].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[346].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[347].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[348].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[349].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[350].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[351].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[352].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[353].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[354].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[355].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[356].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[357].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[358].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[359].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[360].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[361].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[362].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[363].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[364].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[365].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[366].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[367].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[368].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[369].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[370].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[371].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[372].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[373].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[374].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[375].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[376].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[377].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[378].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[379].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[380].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[381].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[382].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[383].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[384].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[385].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[386].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[387].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[388].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[389].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[390].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[391].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[392].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[393].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[394].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[395].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[396].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[397].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[398].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[399].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[400].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[401].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[402].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[403].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[404].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[405].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[406].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[407].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[408].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[409].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[410].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[411].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[412].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[413].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[414].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[415].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[416].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[417].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[418].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[419].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[420].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[421].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[422].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[423].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[424].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[425].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[426].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[427].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[428].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[429].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[430].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[431].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[432].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[433].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[434].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[435].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[436].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[437].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[438].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[439].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[440].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[441].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[442].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[443].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[444].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[445].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[446].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[447].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[448].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_D.slave[449].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      
      env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      
      env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.disable_check(env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.signal_valid_tvalid_check);
    `endif
    `ifdef TB_CONFIG_2
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.signal_valid_tvalid_check);
    `endif
    `ifdef TB_CONFIG_3
      env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.disable_check(env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.signal_valid_tvalid_check);
    `endif

    root.print_topology();
    `uvm_info("end_of_elaboration_phase", "Exiting...", UVM_LOW)
  endfunction: end_of_elaboration_phase


  /**
   * Calculate the pass or fail status for the test in the final phase method of the
   * test. If a UVM_FATAL or UVM_ERROR message has been generated the
   * test will fail.
   */
  function void final_phase(uvm_phase phase);
    uvm_report_server svr;
    `uvm_info("final_phase", "Entered...",UVM_LOW)

    super.final_phase(phase);

    svr = uvm_report_server::get_server();

    if (svr.get_severity_count(UVM_FATAL) +
        svr.get_severity_count(UVM_ERROR) > 0) 
      `uvm_info("final_phase", "\nTest Status : Failed\n", UVM_LOW)
    else
      `uvm_info("final_phase", "\nTest Status : Passed\n", UVM_LOW)

    `uvm_info("final_phase", "Exiting...", UVM_LOW)
  endfunction: final_phase


  function disable_tready_check();
   `uvm_info("BASE_TEST", "Disabling tready check for invalid scenario ...",UVM_LOW)
    env.pf_vf_mux_system_env_H.master[0].monitor.checks.disable_check(env.pf_vf_mux_system_env_H.master[0].monitor.checks.signal_valid_tready_when_tvalid_high_check);
  endfunction


  function enable_vip_error();
   `uvm_info("BASE_TEST", "ENABLE_VIP_ERR ...",UVM_LOW)
    env.pf_vf_mux_system_env_H.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_H.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_D.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
    `ifdef TB_CONFIG_4
      env.pf_vf_mux_system_env_D.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_D.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      
      env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
      
      
      env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.tvalid_low_when_reset_is_active_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif
    `ifdef TB_CONFIG_2
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif
    `ifdef TB_CONFIG_3
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.tvalid_low_when_reset_is_active_check);
    env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.tvalid_low_when_reset_is_active_check);
    `endif

    env.pf_vf_mux_system_env_H.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_H.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[1].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[2].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[3].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[4].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[5].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[6].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[7].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[8].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[9].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[10].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[11].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[12].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[13].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[14].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_D.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[15].monitor.checks.signal_valid_tvalid_check);
    `ifdef TB_CONFIG_4
   env.pf_vf_mux_system_env_D.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[16].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[17].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[18].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[19].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[20].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[21].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[22].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[23].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[24].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[25].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[26].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[27].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[28].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[29].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[30].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[31].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[32].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[33].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[34].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[35].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[36].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[37].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[38].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[39].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[40].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[41].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[42].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[43].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[44].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[45].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[46].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[47].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[48].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[49].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[50].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[51].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[52].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[53].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[54].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[55].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[56].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[57].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[58].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[59].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[60].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[61].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[62].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[63].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[64].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[65].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[66].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[67].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[68].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[69].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[70].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[71].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[72].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[73].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[74].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[75].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[76].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[77].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[78].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[79].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[80].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[81].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[82].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[83].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[84].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[85].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[86].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[87].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[88].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[89].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[90].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[91].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[92].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[93].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[94].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[95].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[96].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[97].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[98].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[99].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[100].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[101].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[102].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[103].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[104].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[105].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[106].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[107].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[108].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[109].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[110].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[111].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[112].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[113].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[114].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[115].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[116].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[117].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[118].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[119].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[120].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[121].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[122].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[123].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[124].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[125].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[126].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[127].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[128].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[129].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[130].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[131].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[132].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[133].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[134].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[135].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[136].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[137].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[138].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[139].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[140].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[141].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[142].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[143].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[144].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[145].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[146].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[147].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[148].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[149].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[150].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[151].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[152].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[153].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[154].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[155].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[156].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[157].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[158].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[159].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[160].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[161].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[162].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[163].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[164].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[165].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[166].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[167].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[168].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[169].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[170].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[171].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[172].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[173].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[174].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[175].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[176].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[177].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[178].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[179].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[180].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[181].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[182].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[183].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[184].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[185].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[186].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[187].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[188].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[189].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[190].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[191].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[192].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[193].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[194].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[195].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[196].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[197].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[198].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[199].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[200].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[201].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[202].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[203].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[204].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[205].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[206].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[207].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[208].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[209].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[210].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[211].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[212].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[213].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[214].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[215].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[216].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[217].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[218].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[219].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[220].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[221].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[222].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[223].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[224].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[225].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[226].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[227].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[228].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[229].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[230].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[231].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[232].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[233].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[234].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[235].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[236].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[237].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[238].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[239].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[240].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[241].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[242].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[243].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[244].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[245].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[246].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[247].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[248].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[249].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[250].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[251].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[252].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[253].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[254].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[255].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[256].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[257].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[258].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[259].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[260].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[261].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[262].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[263].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[264].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[265].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[266].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[267].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[268].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[269].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[270].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[271].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[272].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[273].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[274].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[275].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[276].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[277].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[278].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[279].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[280].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[281].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[282].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[283].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[284].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[285].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[286].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[287].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[288].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[289].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[290].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[291].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[292].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[293].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[294].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[295].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[296].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[297].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[298].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[299].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[300].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[301].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[302].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[303].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[304].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[305].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[306].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[307].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[308].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[309].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[310].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[311].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[312].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[313].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[314].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[315].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[316].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[317].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[318].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[319].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[320].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[321].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[322].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[323].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[324].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[325].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[326].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[327].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[328].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[329].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[330].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[331].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[332].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[333].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[334].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[335].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[336].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[337].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[338].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[339].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[340].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[341].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[342].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[343].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[344].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[345].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[346].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[347].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[348].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[349].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[350].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[351].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[352].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[353].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[354].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[355].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[356].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[357].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[358].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[359].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[360].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[361].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[362].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[363].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[364].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[365].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[366].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[367].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[368].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[369].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[370].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[371].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[372].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[373].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[374].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[375].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[376].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[377].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[378].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[379].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[380].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[381].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[382].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[383].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[384].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[385].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[386].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[387].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[388].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[389].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[390].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[391].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[392].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[393].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[394].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[395].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[396].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[397].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[398].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[399].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[400].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[401].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[402].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[403].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[404].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[405].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[406].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[407].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[408].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[409].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[410].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[411].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[412].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[413].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[414].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[415].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[416].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[417].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[418].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[419].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[420].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[421].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[422].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[423].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[424].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[425].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[426].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[427].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[428].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[429].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[430].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[431].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[432].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[433].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[434].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[435].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[436].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[437].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[438].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[439].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[440].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[441].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[442].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[443].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[444].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[445].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[446].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[447].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[448].monitor.checks.signal_valid_tvalid_check);
   env.pf_vf_mux_system_env_D.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_D.slave[449].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D0.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D1.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      
      env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D2.slave[449].monitor.checks.signal_valid_tvalid_check);
      
      
      env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[0].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[1].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[2].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[3].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[4].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[5].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[6].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[7].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[8].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[9].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[10].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[11].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[12].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[13].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[14].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[15].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[16].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[17].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[18].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[19].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[20].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[21].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[22].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[23].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[24].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[25].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[26].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[27].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[28].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[29].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[30].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[31].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[32].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[33].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[34].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[35].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[36].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[37].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[38].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[39].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[40].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[41].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[42].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[43].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[44].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[45].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[46].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[47].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[48].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[49].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[50].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[51].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[52].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[53].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[54].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[55].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[56].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[57].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[58].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[59].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[60].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[61].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[62].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[63].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[64].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[65].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[66].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[67].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[68].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[69].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[70].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[71].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[72].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[73].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[74].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[75].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[76].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[77].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[78].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[79].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[80].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[81].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[82].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[83].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[84].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[85].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[86].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[87].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[88].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[89].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[90].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[91].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[92].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[93].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[94].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[95].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[96].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[97].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[98].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[99].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[100].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[101].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[102].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[103].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[104].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[105].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[106].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[107].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[108].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[109].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[110].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[111].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[112].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[113].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[114].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[115].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[116].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[117].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[118].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[119].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[120].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[121].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[122].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[123].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[124].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[125].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[126].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[127].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[128].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[129].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[130].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[131].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[132].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[133].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[134].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[135].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[136].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[137].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[138].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[139].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[140].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[141].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[142].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[143].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[144].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[145].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[146].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[147].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[148].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[149].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[150].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[151].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[152].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[153].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[154].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[155].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[156].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[157].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[158].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[159].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[160].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[161].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[162].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[163].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[164].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[165].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[166].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[167].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[168].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[169].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[170].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[171].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[172].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[173].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[174].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[175].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[176].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[177].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[178].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[179].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[180].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[181].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[182].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[183].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[184].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[185].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[186].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[187].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[188].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[189].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[190].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[191].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[192].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[193].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[194].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[195].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[196].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[197].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[198].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[199].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[200].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[201].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[202].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[203].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[204].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[205].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[206].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[207].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[208].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[209].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[210].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[211].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[212].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[213].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[214].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[215].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[216].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[217].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[218].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[219].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[220].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[221].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[222].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[223].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[224].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[225].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[226].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[227].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[228].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[229].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[230].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[231].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[232].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[233].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[234].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[235].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[236].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[237].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[238].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[239].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[240].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[241].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[242].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[243].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[244].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[245].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[246].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[247].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[248].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[249].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[250].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[251].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[252].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[253].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[254].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[255].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[256].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[257].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[258].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[259].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[260].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[261].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[262].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[263].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[264].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[265].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[266].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[267].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[268].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[269].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[270].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[271].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[272].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[273].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[274].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[275].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[276].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[277].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[278].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[279].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[280].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[281].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[282].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[283].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[284].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[285].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[286].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[287].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[288].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[289].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[290].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[291].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[292].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[293].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[294].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[295].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[296].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[297].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[298].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[299].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[300].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[301].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[302].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[303].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[304].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[305].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[306].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[307].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[308].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[309].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[310].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[311].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[312].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[313].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[314].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[315].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[316].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[317].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[318].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[319].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[320].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[321].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[322].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[323].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[324].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[325].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[326].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[327].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[328].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[329].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[330].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[331].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[332].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[333].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[334].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[335].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[336].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[337].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[338].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[339].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[340].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[341].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[342].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[343].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[344].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[345].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[346].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[347].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[348].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[349].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[350].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[351].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[352].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[353].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[354].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[355].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[356].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[357].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[358].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[359].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[360].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[361].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[362].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[363].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[364].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[365].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[366].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[367].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[368].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[369].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[370].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[371].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[372].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[373].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[374].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[375].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[376].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[377].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[378].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[379].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[380].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[381].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[382].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[383].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[384].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[385].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[386].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[387].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[388].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[389].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[390].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[391].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[392].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[393].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[394].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[395].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[396].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[397].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[398].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[399].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[400].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[401].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[402].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[403].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[404].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[405].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[406].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[407].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[408].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[409].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[410].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[411].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[412].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[413].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[414].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[415].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[416].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[417].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[418].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[419].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[420].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[421].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[422].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[423].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[424].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[425].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[426].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[427].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[428].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[429].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[430].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[431].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[432].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[433].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[434].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[435].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[436].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[437].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[438].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[439].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[440].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[441].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[442].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[443].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[444].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[445].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[446].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[447].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[448].monitor.checks.signal_valid_tvalid_check);
      env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.enable_check(env.pf_vf_mux_system_env_TB4_D3.slave[449].monitor.checks.signal_valid_tvalid_check);
   `endif   
    `ifdef TB_CONFIG_2
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.signal_valid_tvalid_check);
    `endif
    `ifdef TB_CONFIG_3
    env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[0].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[1].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[2].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[3].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[4].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[5].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[6].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[7].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[8].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[9].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[10].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[11].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[12].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[13].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[14].monitor.checks.signal_valid_tvalid_check);
    env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.enable_check(env.pf_vf_mux_system_env_DN.slave[15].monitor.checks.signal_valid_tvalid_check);
    `endif

  endfunction

  function final_packet_count_check();
      uvm_config_db#(int)::get(null, "", "no_of_trans", packet_count);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_0.packet_count,0);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1.packet_count,1);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2.packet_count,2);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_3.packet_count,3);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_4.packet_count,4);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_5.packet_count,5);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_6.packet_count,6);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_7.packet_count,7);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_8.packet_count,8);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_9.packet_count,9);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_10.packet_count,10);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_11.packet_count,11);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_12.packet_count,12);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_13.packet_count,13);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_14.packet_count,14);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_15.packet_count,15);
      `ifdef TB_CONFIG_2
        packet_count_check(packet_count,env.pf_vf_mux_scbd_16.packet_count,16);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_17.packet_count,17);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_18.packet_count,18);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_19.packet_count,19);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_20.packet_count,20);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_21.packet_count,21);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_22.packet_count,22);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_23.packet_count,23);
      `elsif TB_CONFIG_3  
        packet_count_check(packet_count,env.pf_vf_mux_scbd_16.packet_count,16);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_17.packet_count,17);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_18.packet_count,18);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_19.packet_count,19);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_20.packet_count,20);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_21.packet_count,21);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_22.packet_count,22);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_23.packet_count,23);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_24.packet_count,24);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_25.packet_count,25);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_26.packet_count,26);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_27.packet_count,27);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_28.packet_count,28);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_29.packet_count,29);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_30.packet_count,30);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_31.packet_count,31);
      `elsif TB_CONFIG_4  
        packet_count_check(packet_count,env.pf_vf_mux_scbd_16.packet_count,16);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_17.packet_count,17);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_18.packet_count,18);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_19.packet_count,19);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_20.packet_count,20);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_21.packet_count,21);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_22.packet_count,22);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_23.packet_count,23);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_24.packet_count,24);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_25.packet_count,25);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_26.packet_count,26);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_27.packet_count,27);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_28.packet_count,28);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_29.packet_count,29);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_30.packet_count,30);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_31.packet_count,31);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_32.packet_count,32);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_33.packet_count,33);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_34.packet_count,34);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_35.packet_count,35);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_36.packet_count,36);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_37.packet_count,37);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_38.packet_count,38);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_39.packet_count,39);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_40.packet_count,40);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_41.packet_count,41);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_42.packet_count,42);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_43.packet_count,43);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_44.packet_count,44);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_45.packet_count,45);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_46.packet_count,46);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_47.packet_count,47);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_48.packet_count,48);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_49.packet_count,49);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_50.packet_count,50);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_51.packet_count,51);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_52.packet_count,52);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_53.packet_count,53);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_54.packet_count,54);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_55.packet_count,55);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_56.packet_count,56);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_57.packet_count,57);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_58.packet_count,58);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_59.packet_count,59);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_60.packet_count,60);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_61.packet_count,61);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_62.packet_count,62);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_63.packet_count,63);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_64.packet_count,64);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_65.packet_count,65);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_66.packet_count,66);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_67.packet_count,67);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_68.packet_count,68);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_69.packet_count,69);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_70.packet_count,70);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_71.packet_count,71);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_72.packet_count,72);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_73.packet_count,73);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_74.packet_count,74);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_75.packet_count,75);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_76.packet_count,76);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_77.packet_count,77);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_78.packet_count,78);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_79.packet_count,79);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_80.packet_count,80);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_81.packet_count,81);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_82.packet_count,82);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_83.packet_count,83);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_84.packet_count,84);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_85.packet_count,85);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_86.packet_count,86);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_87.packet_count,87);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_88.packet_count,88);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_89.packet_count,89);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_90.packet_count,90);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_91.packet_count,91);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_92.packet_count,92);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_93.packet_count,93);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_94.packet_count,94);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_95.packet_count,95);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_96.packet_count,96);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_97.packet_count,97);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_98.packet_count,98);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_99.packet_count,99);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_100.packet_count,100);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_101.packet_count,101);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_102.packet_count,102);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_103.packet_count,103);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_104.packet_count,104);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_105.packet_count,105);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_106.packet_count,106);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_107.packet_count,107);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_108.packet_count,108);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_109.packet_count,109);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_110.packet_count,110);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_111.packet_count,111);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_112.packet_count,112);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_113.packet_count,113);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_114.packet_count,114);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_115.packet_count,115);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_116.packet_count,116);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_117.packet_count,117);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_118.packet_count,118);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_119.packet_count,119);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_120.packet_count,120);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_121.packet_count,121);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_122.packet_count,122);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_123.packet_count,123);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_124.packet_count,124);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_125.packet_count,125);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_126.packet_count,126);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_127.packet_count,127);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_128.packet_count,128);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_129.packet_count,129);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_130.packet_count,130);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_131.packet_count,131);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_132.packet_count,132);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_133.packet_count,133);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_134.packet_count,134);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_135.packet_count,135);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_136.packet_count,136);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_137.packet_count,137);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_138.packet_count,138);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_139.packet_count,139);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_140.packet_count,140);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_141.packet_count,141);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_142.packet_count,142);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_143.packet_count,143);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_144.packet_count,144);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_145.packet_count,145);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_146.packet_count,146);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_147.packet_count,147);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_148.packet_count,148);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_149.packet_count,149);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_150.packet_count,150);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_151.packet_count,151);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_152.packet_count,152);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_153.packet_count,153);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_154.packet_count,154);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_155.packet_count,155);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_156.packet_count,156);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_157.packet_count,157);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_158.packet_count,158);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_159.packet_count,159);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_160.packet_count,160);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_161.packet_count,161);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_162.packet_count,162);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_163.packet_count,163);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_164.packet_count,164);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_165.packet_count,165);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_166.packet_count,166);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_167.packet_count,167);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_168.packet_count,168);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_169.packet_count,169);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_170.packet_count,170);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_171.packet_count,171);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_172.packet_count,172);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_173.packet_count,173);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_174.packet_count,174);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_175.packet_count,175);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_176.packet_count,176);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_177.packet_count,177);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_178.packet_count,178);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_179.packet_count,179);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_180.packet_count,180);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_181.packet_count,181);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_182.packet_count,182);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_183.packet_count,183);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_184.packet_count,184);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_185.packet_count,185);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_186.packet_count,186);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_187.packet_count,187);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_188.packet_count,188);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_189.packet_count,189);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_190.packet_count,190);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_191.packet_count,191);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_192.packet_count,192);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_193.packet_count,193);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_194.packet_count,194);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_195.packet_count,195);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_196.packet_count,196);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_197.packet_count,197);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_198.packet_count,198);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_199.packet_count,199);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_200.packet_count,200);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_201.packet_count,201);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_202.packet_count,202);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_203.packet_count,203);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_204.packet_count,204);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_205.packet_count,205);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_206.packet_count,206);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_207.packet_count,207);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_208.packet_count,208);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_209.packet_count,209);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_210.packet_count,210);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_211.packet_count,211);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_212.packet_count,212);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_213.packet_count,213);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_214.packet_count,214);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_215.packet_count,215);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_216.packet_count,216);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_217.packet_count,217);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_218.packet_count,218);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_219.packet_count,219);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_220.packet_count,220);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_221.packet_count,221);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_222.packet_count,222);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_223.packet_count,223);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_224.packet_count,224);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_225.packet_count,225);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_226.packet_count,226);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_227.packet_count,227);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_228.packet_count,228);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_229.packet_count,229);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_230.packet_count,230);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_231.packet_count,231);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_232.packet_count,232);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_233.packet_count,233);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_234.packet_count,234);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_235.packet_count,235);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_236.packet_count,236);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_237.packet_count,237);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_238.packet_count,238);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_239.packet_count,239);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_240.packet_count,240);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_241.packet_count,241);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_242.packet_count,242);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_243.packet_count,243);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_244.packet_count,244);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_245.packet_count,245);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_246.packet_count,246);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_247.packet_count,247);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_248.packet_count,248);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_249.packet_count,249);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_250.packet_count,250);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_251.packet_count,251);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_252.packet_count,252);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_253.packet_count,253);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_254.packet_count,254);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_255.packet_count,255);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_256.packet_count,256);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_257.packet_count,257);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_258.packet_count,258);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_259.packet_count,259);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_260.packet_count,260);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_261.packet_count,261);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_262.packet_count,262);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_263.packet_count,263);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_264.packet_count,264);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_265.packet_count,265);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_266.packet_count,266);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_267.packet_count,267);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_268.packet_count,268);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_269.packet_count,269);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_270.packet_count,270);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_271.packet_count,271);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_272.packet_count,272);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_273.packet_count,273);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_274.packet_count,274);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_275.packet_count,275);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_276.packet_count,276);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_277.packet_count,277);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_278.packet_count,278);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_279.packet_count,279);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_280.packet_count,280);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_281.packet_count,281);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_282.packet_count,282);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_283.packet_count,283);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_284.packet_count,284);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_285.packet_count,285);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_286.packet_count,286);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_287.packet_count,287);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_288.packet_count,288);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_289.packet_count,289);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_290.packet_count,290);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_291.packet_count,291);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_292.packet_count,292);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_293.packet_count,293);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_294.packet_count,294);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_295.packet_count,295);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_296.packet_count,296);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_297.packet_count,297);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_298.packet_count,298);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_299.packet_count,299);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_300.packet_count,300);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_301.packet_count,301);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_302.packet_count,302);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_303.packet_count,303);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_304.packet_count,304);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_305.packet_count,305);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_306.packet_count,306);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_307.packet_count,307);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_308.packet_count,308);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_309.packet_count,309);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_310.packet_count,310);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_311.packet_count,311);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_312.packet_count,312);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_313.packet_count,313);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_314.packet_count,314);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_315.packet_count,315);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_316.packet_count,316);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_317.packet_count,317);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_318.packet_count,318);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_319.packet_count,319);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_320.packet_count,320);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_321.packet_count,321);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_322.packet_count,322);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_323.packet_count,323);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_324.packet_count,324);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_325.packet_count,325);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_326.packet_count,326);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_327.packet_count,327);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_328.packet_count,328);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_329.packet_count,329);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_330.packet_count,330);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_331.packet_count,331);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_332.packet_count,332);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_333.packet_count,333);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_334.packet_count,334);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_335.packet_count,335);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_336.packet_count,336);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_337.packet_count,337);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_338.packet_count,338);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_339.packet_count,339);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_340.packet_count,340);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_341.packet_count,341);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_342.packet_count,342);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_343.packet_count,343);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_344.packet_count,344);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_345.packet_count,345);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_346.packet_count,346);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_347.packet_count,347);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_348.packet_count,348);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_349.packet_count,349);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_350.packet_count,350);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_351.packet_count,351);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_352.packet_count,352);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_353.packet_count,353);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_354.packet_count,354);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_355.packet_count,355);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_356.packet_count,356);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_357.packet_count,357);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_358.packet_count,358);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_359.packet_count,359);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_360.packet_count,360);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_361.packet_count,361);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_362.packet_count,362);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_363.packet_count,363);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_364.packet_count,364);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_365.packet_count,365);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_366.packet_count,366);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_367.packet_count,367);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_368.packet_count,368);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_369.packet_count,369);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_370.packet_count,370);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_371.packet_count,371);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_372.packet_count,372);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_373.packet_count,373);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_374.packet_count,374);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_375.packet_count,375);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_376.packet_count,376);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_377.packet_count,377);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_378.packet_count,378);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_379.packet_count,379);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_380.packet_count,380);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_381.packet_count,381);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_382.packet_count,382);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_383.packet_count,383);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_384.packet_count,384);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_385.packet_count,385);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_386.packet_count,386);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_387.packet_count,387);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_388.packet_count,388);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_389.packet_count,389);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_390.packet_count,390);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_391.packet_count,391);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_392.packet_count,392);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_393.packet_count,393);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_394.packet_count,394);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_395.packet_count,395);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_396.packet_count,396);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_397.packet_count,397);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_398.packet_count,398);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_399.packet_count,399);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_400.packet_count,400);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_401.packet_count,401);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_402.packet_count,402);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_403.packet_count,403);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_404.packet_count,404);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_405.packet_count,405);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_406.packet_count,406);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_407.packet_count,407);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_408.packet_count,408);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_409.packet_count,409);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_410.packet_count,410);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_411.packet_count,411);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_412.packet_count,412);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_413.packet_count,413);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_414.packet_count,414);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_415.packet_count,415);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_416.packet_count,416);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_417.packet_count,417);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_418.packet_count,418);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_419.packet_count,419);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_420.packet_count,420);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_421.packet_count,421);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_422.packet_count,422);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_423.packet_count,423);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_424.packet_count,424);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_425.packet_count,425);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_426.packet_count,426);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_427.packet_count,427);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_428.packet_count,428);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_429.packet_count,429);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_430.packet_count,430);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_431.packet_count,431);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_432.packet_count,432);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_433.packet_count,433);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_434.packet_count,434);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_435.packet_count,435);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_436.packet_count,436);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_437.packet_count,437);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_438.packet_count,438);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_439.packet_count,439);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_440.packet_count,440);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_441.packet_count,441);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_442.packet_count,442);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_443.packet_count,443);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_444.packet_count,444);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_445.packet_count,445);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_446.packet_count,446);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_447.packet_count,447);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_448.packet_count,448);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_449.packet_count,449);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_450.packet_count,450);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_451.packet_count,451);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_452.packet_count,452);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_453.packet_count,453);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_454.packet_count,454);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_455.packet_count,455);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_456.packet_count,456);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_457.packet_count,457);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_458.packet_count,458);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_459.packet_count,459);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_460.packet_count,460);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_461.packet_count,461);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_462.packet_count,462);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_463.packet_count,463);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_464.packet_count,464);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_465.packet_count,465);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_466.packet_count,466);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_467.packet_count,467);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_468.packet_count,468);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_469.packet_count,469);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_470.packet_count,470);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_471.packet_count,471);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_472.packet_count,472);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_473.packet_count,473);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_474.packet_count,474);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_475.packet_count,475);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_476.packet_count,476);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_477.packet_count,477);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_478.packet_count,478);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_479.packet_count,479);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_480.packet_count,480);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_481.packet_count,481);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_482.packet_count,482);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_483.packet_count,483);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_484.packet_count,484);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_485.packet_count,485);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_486.packet_count,486);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_487.packet_count,487);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_488.packet_count,488);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_489.packet_count,489);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_490.packet_count,490);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_491.packet_count,491);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_492.packet_count,492);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_493.packet_count,493);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_494.packet_count,494);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_495.packet_count,495);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_496.packet_count,496);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_497.packet_count,497);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_498.packet_count,498);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_499.packet_count,499);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_500.packet_count,500);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_501.packet_count,501);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_502.packet_count,502);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_503.packet_count,503);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_504.packet_count,504);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_505.packet_count,505);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_506.packet_count,506);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_507.packet_count,507);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_508.packet_count,508);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_509.packet_count,509);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_510.packet_count,510);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_511.packet_count,511);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_512.packet_count,512);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_513.packet_count,513);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_514.packet_count,514);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_515.packet_count,515);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_516.packet_count,516);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_517.packet_count,517);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_518.packet_count,518);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_519.packet_count,519);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_520.packet_count,520);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_521.packet_count,521);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_522.packet_count,522);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_523.packet_count,523);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_524.packet_count,524);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_525.packet_count,525);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_526.packet_count,526);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_527.packet_count,527);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_528.packet_count,528);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_529.packet_count,529);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_530.packet_count,530);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_531.packet_count,531);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_532.packet_count,532);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_533.packet_count,533);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_534.packet_count,534);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_535.packet_count,535);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_536.packet_count,536);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_537.packet_count,537);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_538.packet_count,538);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_539.packet_count,539);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_540.packet_count,540);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_541.packet_count,541);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_542.packet_count,542);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_543.packet_count,543);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_544.packet_count,544);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_545.packet_count,545);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_546.packet_count,546);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_547.packet_count,547);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_548.packet_count,548);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_549.packet_count,549);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_550.packet_count,550);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_551.packet_count,551);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_552.packet_count,552);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_553.packet_count,553);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_554.packet_count,554);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_555.packet_count,555);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_556.packet_count,556);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_557.packet_count,557);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_558.packet_count,558);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_559.packet_count,559);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_560.packet_count,560);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_561.packet_count,561);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_562.packet_count,562);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_563.packet_count,563);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_564.packet_count,564);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_565.packet_count,565);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_566.packet_count,566);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_567.packet_count,567);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_568.packet_count,568);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_569.packet_count,569);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_570.packet_count,570);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_571.packet_count,571);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_572.packet_count,572);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_573.packet_count,573);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_574.packet_count,574);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_575.packet_count,575);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_576.packet_count,576);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_577.packet_count,577);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_578.packet_count,578);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_579.packet_count,579);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_580.packet_count,580);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_581.packet_count,581);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_582.packet_count,582);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_583.packet_count,583);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_584.packet_count,584);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_585.packet_count,585);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_586.packet_count,586);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_587.packet_count,587);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_588.packet_count,588);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_589.packet_count,589);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_590.packet_count,590);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_591.packet_count,591);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_592.packet_count,592);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_593.packet_count,593);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_594.packet_count,594);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_595.packet_count,595);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_596.packet_count,596);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_597.packet_count,597);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_598.packet_count,598);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_599.packet_count,599);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_600.packet_count,600);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_601.packet_count,601);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_602.packet_count,602);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_603.packet_count,603);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_604.packet_count,604);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_605.packet_count,605);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_606.packet_count,606);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_607.packet_count,607);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_608.packet_count,608);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_609.packet_count,609);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_610.packet_count,610);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_611.packet_count,611);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_612.packet_count,612);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_613.packet_count,613);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_614.packet_count,614);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_615.packet_count,615);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_616.packet_count,616);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_617.packet_count,617);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_618.packet_count,618);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_619.packet_count,619);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_620.packet_count,620);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_621.packet_count,621);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_622.packet_count,622);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_623.packet_count,623);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_624.packet_count,624);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_625.packet_count,625);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_626.packet_count,626);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_627.packet_count,627);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_628.packet_count,628);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_629.packet_count,629);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_630.packet_count,630);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_631.packet_count,631);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_632.packet_count,632);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_633.packet_count,633);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_634.packet_count,634);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_635.packet_count,635);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_636.packet_count,636);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_637.packet_count,637);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_638.packet_count,638);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_639.packet_count,639);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_640.packet_count,640);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_641.packet_count,641);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_642.packet_count,642);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_643.packet_count,643);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_644.packet_count,644);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_645.packet_count,645);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_646.packet_count,646);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_647.packet_count,647);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_648.packet_count,648);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_649.packet_count,649);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_650.packet_count,650);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_651.packet_count,651);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_652.packet_count,652);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_653.packet_count,653);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_654.packet_count,654);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_655.packet_count,655);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_656.packet_count,656);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_657.packet_count,657);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_658.packet_count,658);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_659.packet_count,659);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_660.packet_count,660);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_661.packet_count,661);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_662.packet_count,662);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_663.packet_count,663);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_664.packet_count,664);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_665.packet_count,665);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_666.packet_count,666);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_667.packet_count,667);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_668.packet_count,668);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_669.packet_count,669);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_670.packet_count,670);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_671.packet_count,671);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_672.packet_count,672);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_673.packet_count,673);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_674.packet_count,674);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_675.packet_count,675);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_676.packet_count,676);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_677.packet_count,677);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_678.packet_count,678);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_679.packet_count,679);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_680.packet_count,680);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_681.packet_count,681);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_682.packet_count,682);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_683.packet_count,683);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_684.packet_count,684);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_685.packet_count,685);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_686.packet_count,686);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_687.packet_count,687);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_688.packet_count,688);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_689.packet_count,689);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_690.packet_count,690);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_691.packet_count,691);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_692.packet_count,692);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_693.packet_count,693);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_694.packet_count,694);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_695.packet_count,695);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_696.packet_count,696);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_697.packet_count,697);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_698.packet_count,698);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_699.packet_count,699);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_700.packet_count,700);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_701.packet_count,701);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_702.packet_count,702);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_703.packet_count,703);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_704.packet_count,704);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_705.packet_count,705);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_706.packet_count,706);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_707.packet_count,707);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_708.packet_count,708);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_709.packet_count,709);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_710.packet_count,710);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_711.packet_count,711);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_712.packet_count,712);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_713.packet_count,713);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_714.packet_count,714);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_715.packet_count,715);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_716.packet_count,716);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_717.packet_count,717);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_718.packet_count,718);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_719.packet_count,719);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_720.packet_count,720);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_721.packet_count,721);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_722.packet_count,722);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_723.packet_count,723);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_724.packet_count,724);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_725.packet_count,725);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_726.packet_count,726);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_727.packet_count,727);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_728.packet_count,728);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_729.packet_count,729);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_730.packet_count,730);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_731.packet_count,731);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_732.packet_count,732);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_733.packet_count,733);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_734.packet_count,734);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_735.packet_count,735);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_736.packet_count,736);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_737.packet_count,737);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_738.packet_count,738);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_739.packet_count,739);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_740.packet_count,740);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_741.packet_count,741);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_742.packet_count,742);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_743.packet_count,743);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_744.packet_count,744);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_745.packet_count,745);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_746.packet_count,746);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_747.packet_count,747);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_748.packet_count,748);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_749.packet_count,749);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_750.packet_count,750);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_751.packet_count,751);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_752.packet_count,752);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_753.packet_count,753);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_754.packet_count,754);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_755.packet_count,755);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_756.packet_count,756);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_757.packet_count,757);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_758.packet_count,758);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_759.packet_count,759);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_760.packet_count,760);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_761.packet_count,761);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_762.packet_count,762);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_763.packet_count,763);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_764.packet_count,764);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_765.packet_count,765);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_766.packet_count,766);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_767.packet_count,767);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_768.packet_count,768);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_769.packet_count,769);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_770.packet_count,770);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_771.packet_count,771);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_772.packet_count,772);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_773.packet_count,773);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_774.packet_count,774);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_775.packet_count,775);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_776.packet_count,776);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_777.packet_count,777);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_778.packet_count,778);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_779.packet_count,779);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_780.packet_count,780);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_781.packet_count,781);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_782.packet_count,782);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_783.packet_count,783);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_784.packet_count,784);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_785.packet_count,785);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_786.packet_count,786);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_787.packet_count,787);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_788.packet_count,788);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_789.packet_count,789);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_790.packet_count,790);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_791.packet_count,791);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_792.packet_count,792);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_793.packet_count,793);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_794.packet_count,794);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_795.packet_count,795);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_796.packet_count,796);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_797.packet_count,797);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_798.packet_count,798);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_799.packet_count,799);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_800.packet_count,800);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_801.packet_count,801);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_802.packet_count,802);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_803.packet_count,803);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_804.packet_count,804);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_805.packet_count,805);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_806.packet_count,806);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_807.packet_count,807);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_808.packet_count,808);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_809.packet_count,809);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_810.packet_count,810);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_811.packet_count,811);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_812.packet_count,812);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_813.packet_count,813);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_814.packet_count,814);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_815.packet_count,815);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_816.packet_count,816);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_817.packet_count,817);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_818.packet_count,818);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_819.packet_count,819);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_820.packet_count,820);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_821.packet_count,821);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_822.packet_count,822);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_823.packet_count,823);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_824.packet_count,824);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_825.packet_count,825);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_826.packet_count,826);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_827.packet_count,827);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_828.packet_count,828);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_829.packet_count,829);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_830.packet_count,830);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_831.packet_count,831);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_832.packet_count,832);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_833.packet_count,833);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_834.packet_count,834);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_835.packet_count,835);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_836.packet_count,836);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_837.packet_count,837);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_838.packet_count,838);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_839.packet_count,839);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_840.packet_count,840);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_841.packet_count,841);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_842.packet_count,842);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_843.packet_count,843);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_844.packet_count,844);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_845.packet_count,845);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_846.packet_count,846);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_847.packet_count,847);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_848.packet_count,848);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_849.packet_count,849);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_850.packet_count,850);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_851.packet_count,851);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_852.packet_count,852);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_853.packet_count,853);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_854.packet_count,854);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_855.packet_count,855);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_856.packet_count,856);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_857.packet_count,857);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_858.packet_count,858);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_859.packet_count,859);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_860.packet_count,860);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_861.packet_count,861);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_862.packet_count,862);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_863.packet_count,863);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_864.packet_count,864);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_865.packet_count,865);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_866.packet_count,866);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_867.packet_count,867);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_868.packet_count,868);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_869.packet_count,869);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_870.packet_count,870);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_871.packet_count,871);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_872.packet_count,872);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_873.packet_count,873);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_874.packet_count,874);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_875.packet_count,875);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_876.packet_count,876);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_877.packet_count,877);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_878.packet_count,878);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_879.packet_count,879);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_880.packet_count,880);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_881.packet_count,881);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_882.packet_count,882);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_883.packet_count,883);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_884.packet_count,884);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_885.packet_count,885);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_886.packet_count,886);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_887.packet_count,887);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_888.packet_count,888);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_889.packet_count,889);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_890.packet_count,890);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_891.packet_count,891);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_892.packet_count,892);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_893.packet_count,893);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_894.packet_count,894);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_895.packet_count,895);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_896.packet_count,896);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_897.packet_count,897);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_898.packet_count,898);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_899.packet_count,899);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_900.packet_count,900);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_901.packet_count,901);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_902.packet_count,902);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_903.packet_count,903);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_904.packet_count,904);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_905.packet_count,905);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_906.packet_count,906);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_907.packet_count,907);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_908.packet_count,908);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_909.packet_count,909);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_910.packet_count,910);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_911.packet_count,911);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_912.packet_count,912);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_913.packet_count,913);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_914.packet_count,914);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_915.packet_count,915);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_916.packet_count,916);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_917.packet_count,917);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_918.packet_count,918);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_919.packet_count,919);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_920.packet_count,920);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_921.packet_count,921);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_922.packet_count,922);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_923.packet_count,923);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_924.packet_count,924);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_925.packet_count,925);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_926.packet_count,926);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_927.packet_count,927);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_928.packet_count,928);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_929.packet_count,929);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_930.packet_count,930);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_931.packet_count,931);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_932.packet_count,932);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_933.packet_count,933);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_934.packet_count,934);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_935.packet_count,935);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_936.packet_count,936);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_937.packet_count,937);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_938.packet_count,938);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_939.packet_count,939);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_940.packet_count,940);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_941.packet_count,941);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_942.packet_count,942);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_943.packet_count,943);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_944.packet_count,944);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_945.packet_count,945);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_946.packet_count,946);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_947.packet_count,947);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_948.packet_count,948);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_949.packet_count,949);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_950.packet_count,950);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_951.packet_count,951);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_952.packet_count,952);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_953.packet_count,953);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_954.packet_count,954);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_955.packet_count,955);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_956.packet_count,956);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_957.packet_count,957);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_958.packet_count,958);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_959.packet_count,959);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_960.packet_count,960);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_961.packet_count,961);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_962.packet_count,962);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_963.packet_count,963);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_964.packet_count,964);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_965.packet_count,965);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_966.packet_count,966);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_967.packet_count,967);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_968.packet_count,968);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_969.packet_count,969);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_970.packet_count,970);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_971.packet_count,971);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_972.packet_count,972);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_973.packet_count,973);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_974.packet_count,974);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_975.packet_count,975);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_976.packet_count,976);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_977.packet_count,977);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_978.packet_count,978);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_979.packet_count,979);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_980.packet_count,980);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_981.packet_count,981);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_982.packet_count,982);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_983.packet_count,983);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_984.packet_count,984);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_985.packet_count,985);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_986.packet_count,986);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_987.packet_count,987);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_988.packet_count,988);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_989.packet_count,989);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_990.packet_count,990);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_991.packet_count,991);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_992.packet_count,992);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_993.packet_count,993);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_994.packet_count,994);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_995.packet_count,995);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_996.packet_count,996);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_997.packet_count,997);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_998.packet_count,998);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_999.packet_count,999);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1000.packet_count,1000);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1001.packet_count,1001);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1002.packet_count,1002);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1003.packet_count,1003);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1004.packet_count,1004);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1005.packet_count,1005);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1006.packet_count,1006);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1007.packet_count,1007);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1008.packet_count,1008);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1009.packet_count,1009);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1010.packet_count,1010);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1011.packet_count,1011);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1012.packet_count,1012);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1013.packet_count,1013);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1014.packet_count,1014);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1015.packet_count,1015);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1016.packet_count,1016);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1017.packet_count,1017);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1018.packet_count,1018);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1019.packet_count,1019);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1020.packet_count,1020);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1021.packet_count,1021);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1022.packet_count,1022);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1023.packet_count,1023);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1024.packet_count,1024);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1025.packet_count,1025);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1026.packet_count,1026);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1027.packet_count,1027);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1028.packet_count,1028);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1029.packet_count,1029);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1030.packet_count,1030);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1031.packet_count,1031);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1032.packet_count,1032);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1033.packet_count,1033);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1034.packet_count,1034);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1035.packet_count,1035);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1036.packet_count,1036);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1037.packet_count,1037);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1038.packet_count,1038);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1039.packet_count,1039);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1040.packet_count,1040);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1041.packet_count,1041);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1042.packet_count,1042);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1043.packet_count,1043);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1044.packet_count,1044);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1045.packet_count,1045);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1046.packet_count,1046);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1047.packet_count,1047);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1048.packet_count,1048);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1049.packet_count,1049);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1050.packet_count,1050);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1051.packet_count,1051);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1052.packet_count,1052);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1053.packet_count,1053);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1054.packet_count,1054);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1055.packet_count,1055);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1056.packet_count,1056);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1057.packet_count,1057);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1058.packet_count,1058);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1059.packet_count,1059);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1060.packet_count,1060);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1061.packet_count,1061);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1062.packet_count,1062);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1063.packet_count,1063);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1064.packet_count,1064);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1065.packet_count,1065);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1066.packet_count,1066);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1067.packet_count,1067);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1068.packet_count,1068);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1069.packet_count,1069);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1070.packet_count,1070);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1071.packet_count,1071);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1072.packet_count,1072);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1073.packet_count,1073);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1074.packet_count,1074);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1075.packet_count,1075);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1076.packet_count,1076);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1077.packet_count,1077);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1078.packet_count,1078);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1079.packet_count,1079);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1080.packet_count,1080);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1081.packet_count,1081);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1082.packet_count,1082);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1083.packet_count,1083);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1084.packet_count,1084);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1085.packet_count,1085);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1086.packet_count,1086);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1087.packet_count,1087);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1088.packet_count,1088);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1089.packet_count,1089);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1090.packet_count,1090);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1091.packet_count,1091);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1092.packet_count,1092);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1093.packet_count,1093);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1094.packet_count,1094);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1095.packet_count,1095);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1096.packet_count,1096);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1097.packet_count,1097);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1098.packet_count,1098);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1099.packet_count,1099);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1100.packet_count,1100);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1101.packet_count,1101);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1102.packet_count,1102);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1103.packet_count,1103);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1104.packet_count,1104);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1105.packet_count,1105);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1106.packet_count,1106);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1107.packet_count,1107);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1108.packet_count,1108);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1109.packet_count,1109);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1110.packet_count,1110);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1111.packet_count,1111);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1112.packet_count,1112);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1113.packet_count,1113);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1114.packet_count,1114);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1115.packet_count,1115);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1116.packet_count,1116);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1117.packet_count,1117);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1118.packet_count,1118);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1119.packet_count,1119);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1120.packet_count,1120);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1121.packet_count,1121);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1122.packet_count,1122);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1123.packet_count,1123);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1124.packet_count,1124);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1125.packet_count,1125);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1126.packet_count,1126);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1127.packet_count,1127);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1128.packet_count,1128);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1129.packet_count,1129);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1130.packet_count,1130);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1131.packet_count,1131);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1132.packet_count,1132);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1133.packet_count,1133);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1134.packet_count,1134);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1135.packet_count,1135);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1136.packet_count,1136);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1137.packet_count,1137);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1138.packet_count,1138);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1139.packet_count,1139);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1140.packet_count,1140);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1141.packet_count,1141);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1142.packet_count,1142);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1143.packet_count,1143);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1144.packet_count,1144);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1145.packet_count,1145);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1146.packet_count,1146);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1147.packet_count,1147);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1148.packet_count,1148);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1149.packet_count,1149);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1150.packet_count,1150);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1151.packet_count,1151);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1152.packet_count,1152);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1153.packet_count,1153);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1154.packet_count,1154);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1155.packet_count,1155);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1156.packet_count,1156);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1157.packet_count,1157);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1158.packet_count,1158);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1159.packet_count,1159);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1160.packet_count,1160);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1161.packet_count,1161);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1162.packet_count,1162);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1163.packet_count,1163);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1164.packet_count,1164);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1165.packet_count,1165);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1166.packet_count,1166);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1167.packet_count,1167);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1168.packet_count,1168);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1169.packet_count,1169);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1170.packet_count,1170);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1171.packet_count,1171);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1172.packet_count,1172);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1173.packet_count,1173);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1174.packet_count,1174);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1175.packet_count,1175);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1176.packet_count,1176);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1177.packet_count,1177);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1178.packet_count,1178);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1179.packet_count,1179);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1180.packet_count,1180);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1181.packet_count,1181);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1182.packet_count,1182);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1183.packet_count,1183);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1184.packet_count,1184);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1185.packet_count,1185);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1186.packet_count,1186);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1187.packet_count,1187);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1188.packet_count,1188);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1189.packet_count,1189);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1190.packet_count,1190);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1191.packet_count,1191);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1192.packet_count,1192);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1193.packet_count,1193);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1194.packet_count,1194);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1195.packet_count,1195);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1196.packet_count,1196);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1197.packet_count,1197);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1198.packet_count,1198);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1199.packet_count,1199);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1200.packet_count,1200);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1201.packet_count,1201);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1202.packet_count,1202);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1203.packet_count,1203);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1204.packet_count,1204);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1205.packet_count,1205);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1206.packet_count,1206);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1207.packet_count,1207);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1208.packet_count,1208);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1209.packet_count,1209);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1210.packet_count,1210);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1211.packet_count,1211);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1212.packet_count,1212);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1213.packet_count,1213);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1214.packet_count,1214);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1215.packet_count,1215);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1216.packet_count,1216);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1217.packet_count,1217);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1218.packet_count,1218);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1219.packet_count,1219);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1220.packet_count,1220);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1221.packet_count,1221);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1222.packet_count,1222);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1223.packet_count,1223);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1224.packet_count,1224);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1225.packet_count,1225);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1226.packet_count,1226);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1227.packet_count,1227);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1228.packet_count,1228);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1229.packet_count,1229);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1230.packet_count,1230);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1231.packet_count,1231);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1232.packet_count,1232);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1233.packet_count,1233);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1234.packet_count,1234);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1235.packet_count,1235);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1236.packet_count,1236);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1237.packet_count,1237);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1238.packet_count,1238);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1239.packet_count,1239);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1240.packet_count,1240);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1241.packet_count,1241);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1242.packet_count,1242);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1243.packet_count,1243);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1244.packet_count,1244);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1245.packet_count,1245);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1246.packet_count,1246);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1247.packet_count,1247);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1248.packet_count,1248);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1249.packet_count,1249);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1250.packet_count,1250);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1251.packet_count,1251);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1252.packet_count,1252);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1253.packet_count,1253);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1254.packet_count,1254);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1255.packet_count,1255);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1256.packet_count,1256);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1257.packet_count,1257);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1258.packet_count,1258);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1259.packet_count,1259);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1260.packet_count,1260);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1261.packet_count,1261);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1262.packet_count,1262);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1263.packet_count,1263);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1264.packet_count,1264);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1265.packet_count,1265);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1266.packet_count,1266);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1267.packet_count,1267);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1268.packet_count,1268);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1269.packet_count,1269);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1270.packet_count,1270);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1271.packet_count,1271);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1272.packet_count,1272);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1273.packet_count,1273);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1274.packet_count,1274);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1275.packet_count,1275);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1276.packet_count,1276);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1277.packet_count,1277);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1278.packet_count,1278);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1279.packet_count,1279);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1280.packet_count,1280);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1281.packet_count,1281);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1282.packet_count,1282);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1283.packet_count,1283);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1284.packet_count,1284);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1285.packet_count,1285);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1286.packet_count,1286);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1287.packet_count,1287);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1288.packet_count,1288);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1289.packet_count,1289);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1290.packet_count,1290);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1291.packet_count,1291);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1292.packet_count,1292);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1293.packet_count,1293);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1294.packet_count,1294);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1295.packet_count,1295);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1296.packet_count,1296);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1297.packet_count,1297);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1298.packet_count,1298);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1299.packet_count,1299);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1300.packet_count,1300);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1301.packet_count,1301);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1302.packet_count,1302);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1303.packet_count,1303);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1304.packet_count,1304);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1305.packet_count,1305);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1306.packet_count,1306);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1307.packet_count,1307);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1308.packet_count,1308);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1309.packet_count,1309);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1310.packet_count,1310);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1311.packet_count,1311);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1312.packet_count,1312);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1313.packet_count,1313);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1314.packet_count,1314);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1315.packet_count,1315);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1316.packet_count,1316);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1317.packet_count,1317);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1318.packet_count,1318);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1319.packet_count,1319);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1320.packet_count,1320);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1321.packet_count,1321);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1322.packet_count,1322);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1323.packet_count,1323);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1324.packet_count,1324);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1325.packet_count,1325);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1326.packet_count,1326);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1327.packet_count,1327);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1328.packet_count,1328);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1329.packet_count,1329);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1330.packet_count,1330);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1331.packet_count,1331);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1332.packet_count,1332);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1333.packet_count,1333);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1334.packet_count,1334);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1335.packet_count,1335);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1336.packet_count,1336);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1337.packet_count,1337);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1338.packet_count,1338);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1339.packet_count,1339);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1340.packet_count,1340);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1341.packet_count,1341);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1342.packet_count,1342);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1343.packet_count,1343);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1344.packet_count,1344);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1345.packet_count,1345);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1346.packet_count,1346);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1347.packet_count,1347);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1348.packet_count,1348);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1349.packet_count,1349);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1350.packet_count,1350);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1351.packet_count,1351);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1352.packet_count,1352);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1353.packet_count,1353);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1354.packet_count,1354);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1355.packet_count,1355);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1356.packet_count,1356);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1357.packet_count,1357);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1358.packet_count,1358);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1359.packet_count,1359);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1360.packet_count,1360);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1361.packet_count,1361);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1362.packet_count,1362);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1363.packet_count,1363);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1364.packet_count,1364);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1365.packet_count,1365);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1366.packet_count,1366);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1367.packet_count,1367);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1368.packet_count,1368);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1369.packet_count,1369);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1370.packet_count,1370);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1371.packet_count,1371);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1372.packet_count,1372);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1373.packet_count,1373);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1374.packet_count,1374);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1375.packet_count,1375);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1376.packet_count,1376);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1377.packet_count,1377);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1378.packet_count,1378);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1379.packet_count,1379);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1380.packet_count,1380);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1381.packet_count,1381);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1382.packet_count,1382);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1383.packet_count,1383);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1384.packet_count,1384);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1385.packet_count,1385);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1386.packet_count,1386);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1387.packet_count,1387);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1388.packet_count,1388);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1389.packet_count,1389);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1390.packet_count,1390);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1391.packet_count,1391);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1392.packet_count,1392);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1393.packet_count,1393);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1394.packet_count,1394);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1395.packet_count,1395);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1396.packet_count,1396);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1397.packet_count,1397);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1398.packet_count,1398);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1399.packet_count,1399);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1400.packet_count,1400);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1401.packet_count,1401);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1402.packet_count,1402);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1403.packet_count,1403);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1404.packet_count,1404);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1405.packet_count,1405);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1406.packet_count,1406);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1407.packet_count,1407);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1408.packet_count,1408);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1409.packet_count,1409);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1410.packet_count,1410);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1411.packet_count,1411);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1412.packet_count,1412);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1413.packet_count,1413);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1414.packet_count,1414);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1415.packet_count,1415);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1416.packet_count,1416);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1417.packet_count,1417);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1418.packet_count,1418);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1419.packet_count,1419);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1420.packet_count,1420);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1421.packet_count,1421);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1422.packet_count,1422);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1423.packet_count,1423);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1424.packet_count,1424);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1425.packet_count,1425);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1426.packet_count,1426);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1427.packet_count,1427);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1428.packet_count,1428);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1429.packet_count,1429);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1430.packet_count,1430);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1431.packet_count,1431);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1432.packet_count,1432);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1433.packet_count,1433);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1434.packet_count,1434);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1435.packet_count,1435);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1436.packet_count,1436);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1437.packet_count,1437);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1438.packet_count,1438);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1439.packet_count,1439);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1440.packet_count,1440);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1441.packet_count,1441);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1442.packet_count,1442);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1443.packet_count,1443);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1444.packet_count,1444);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1445.packet_count,1445);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1446.packet_count,1446);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1447.packet_count,1447);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1448.packet_count,1448);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1449.packet_count,1449);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1450.packet_count,1450);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1451.packet_count,1451);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1452.packet_count,1452);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1453.packet_count,1453);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1454.packet_count,1454);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1455.packet_count,1455);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1456.packet_count,1456);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1457.packet_count,1457);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1458.packet_count,1458);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1459.packet_count,1459);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1460.packet_count,1460);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1461.packet_count,1461);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1462.packet_count,1462);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1463.packet_count,1463);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1464.packet_count,1464);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1465.packet_count,1465);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1466.packet_count,1466);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1467.packet_count,1467);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1468.packet_count,1468);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1469.packet_count,1469);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1470.packet_count,1470);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1471.packet_count,1471);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1472.packet_count,1472);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1473.packet_count,1473);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1474.packet_count,1474);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1475.packet_count,1475);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1476.packet_count,1476);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1477.packet_count,1477);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1478.packet_count,1478);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1479.packet_count,1479);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1480.packet_count,1480);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1481.packet_count,1481);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1482.packet_count,1482);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1483.packet_count,1483);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1484.packet_count,1484);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1485.packet_count,1485);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1486.packet_count,1486);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1487.packet_count,1487);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1488.packet_count,1488);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1489.packet_count,1489);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1490.packet_count,1490);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1491.packet_count,1491);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1492.packet_count,1492);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1493.packet_count,1493);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1494.packet_count,1494);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1495.packet_count,1495);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1496.packet_count,1496);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1497.packet_count,1497);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1498.packet_count,1498);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1499.packet_count,1499);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1500.packet_count,1500);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1501.packet_count,1501);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1502.packet_count,1502);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1503.packet_count,1503);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1504.packet_count,1504);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1505.packet_count,1505);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1506.packet_count,1506);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1507.packet_count,1507);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1508.packet_count,1508);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1509.packet_count,1509);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1510.packet_count,1510);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1511.packet_count,1511);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1512.packet_count,1512);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1513.packet_count,1513);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1514.packet_count,1514);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1515.packet_count,1515);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1516.packet_count,1516);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1517.packet_count,1517);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1518.packet_count,1518);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1519.packet_count,1519);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1520.packet_count,1520);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1521.packet_count,1521);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1522.packet_count,1522);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1523.packet_count,1523);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1524.packet_count,1524);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1525.packet_count,1525);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1526.packet_count,1526);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1527.packet_count,1527);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1528.packet_count,1528);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1529.packet_count,1529);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1530.packet_count,1530);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1531.packet_count,1531);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1532.packet_count,1532);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1533.packet_count,1533);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1534.packet_count,1534);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1535.packet_count,1535);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1536.packet_count,1536);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1537.packet_count,1537);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1538.packet_count,1538);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1539.packet_count,1539);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1540.packet_count,1540);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1541.packet_count,1541);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1542.packet_count,1542);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1543.packet_count,1543);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1544.packet_count,1544);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1545.packet_count,1545);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1546.packet_count,1546);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1547.packet_count,1547);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1548.packet_count,1548);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1549.packet_count,1549);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1550.packet_count,1550);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1551.packet_count,1551);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1552.packet_count,1552);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1553.packet_count,1553);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1554.packet_count,1554);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1555.packet_count,1555);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1556.packet_count,1556);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1557.packet_count,1557);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1558.packet_count,1558);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1559.packet_count,1559);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1560.packet_count,1560);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1561.packet_count,1561);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1562.packet_count,1562);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1563.packet_count,1563);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1564.packet_count,1564);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1565.packet_count,1565);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1566.packet_count,1566);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1567.packet_count,1567);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1568.packet_count,1568);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1569.packet_count,1569);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1570.packet_count,1570);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1571.packet_count,1571);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1572.packet_count,1572);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1573.packet_count,1573);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1574.packet_count,1574);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1575.packet_count,1575);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1576.packet_count,1576);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1577.packet_count,1577);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1578.packet_count,1578);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1579.packet_count,1579);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1580.packet_count,1580);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1581.packet_count,1581);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1582.packet_count,1582);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1583.packet_count,1583);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1584.packet_count,1584);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1585.packet_count,1585);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1586.packet_count,1586);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1587.packet_count,1587);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1588.packet_count,1588);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1589.packet_count,1589);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1590.packet_count,1590);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1591.packet_count,1591);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1592.packet_count,1592);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1593.packet_count,1593);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1594.packet_count,1594);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1595.packet_count,1595);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1596.packet_count,1596);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1597.packet_count,1597);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1598.packet_count,1598);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1599.packet_count,1599);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1600.packet_count,1600);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1601.packet_count,1601);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1602.packet_count,1602);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1603.packet_count,1603);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1604.packet_count,1604);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1605.packet_count,1605);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1606.packet_count,1606);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1607.packet_count,1607);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1608.packet_count,1608);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1609.packet_count,1609);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1610.packet_count,1610);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1611.packet_count,1611);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1612.packet_count,1612);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1613.packet_count,1613);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1614.packet_count,1614);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1615.packet_count,1615);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1616.packet_count,1616);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1617.packet_count,1617);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1618.packet_count,1618);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1619.packet_count,1619);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1620.packet_count,1620);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1621.packet_count,1621);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1622.packet_count,1622);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1623.packet_count,1623);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1624.packet_count,1624);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1625.packet_count,1625);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1626.packet_count,1626);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1627.packet_count,1627);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1628.packet_count,1628);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1629.packet_count,1629);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1630.packet_count,1630);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1631.packet_count,1631);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1632.packet_count,1632);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1633.packet_count,1633);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1634.packet_count,1634);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1635.packet_count,1635);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1636.packet_count,1636);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1637.packet_count,1637);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1638.packet_count,1638);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1639.packet_count,1639);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1640.packet_count,1640);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1641.packet_count,1641);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1642.packet_count,1642);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1643.packet_count,1643);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1644.packet_count,1644);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1645.packet_count,1645);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1646.packet_count,1646);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1647.packet_count,1647);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1648.packet_count,1648);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1649.packet_count,1649);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1650.packet_count,1650);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1651.packet_count,1651);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1652.packet_count,1652);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1653.packet_count,1653);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1654.packet_count,1654);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1655.packet_count,1655);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1656.packet_count,1656);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1657.packet_count,1657);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1658.packet_count,1658);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1659.packet_count,1659);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1660.packet_count,1660);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1661.packet_count,1661);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1662.packet_count,1662);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1663.packet_count,1663);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1664.packet_count,1664);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1665.packet_count,1665);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1666.packet_count,1666);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1667.packet_count,1667);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1668.packet_count,1668);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1669.packet_count,1669);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1670.packet_count,1670);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1671.packet_count,1671);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1672.packet_count,1672);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1673.packet_count,1673);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1674.packet_count,1674);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1675.packet_count,1675);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1676.packet_count,1676);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1677.packet_count,1677);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1678.packet_count,1678);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1679.packet_count,1679);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1680.packet_count,1680);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1681.packet_count,1681);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1682.packet_count,1682);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1683.packet_count,1683);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1684.packet_count,1684);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1685.packet_count,1685);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1686.packet_count,1686);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1687.packet_count,1687);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1688.packet_count,1688);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1689.packet_count,1689);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1690.packet_count,1690);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1691.packet_count,1691);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1692.packet_count,1692);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1693.packet_count,1693);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1694.packet_count,1694);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1695.packet_count,1695);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1696.packet_count,1696);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1697.packet_count,1697);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1698.packet_count,1698);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1699.packet_count,1699);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1700.packet_count,1700);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1701.packet_count,1701);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1702.packet_count,1702);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1703.packet_count,1703);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1704.packet_count,1704);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1705.packet_count,1705);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1706.packet_count,1706);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1707.packet_count,1707);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1708.packet_count,1708);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1709.packet_count,1709);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1710.packet_count,1710);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1711.packet_count,1711);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1712.packet_count,1712);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1713.packet_count,1713);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1714.packet_count,1714);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1715.packet_count,1715);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1716.packet_count,1716);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1717.packet_count,1717);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1718.packet_count,1718);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1719.packet_count,1719);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1720.packet_count,1720);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1721.packet_count,1721);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1722.packet_count,1722);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1723.packet_count,1723);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1724.packet_count,1724);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1725.packet_count,1725);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1726.packet_count,1726);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1727.packet_count,1727);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1728.packet_count,1728);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1729.packet_count,1729);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1730.packet_count,1730);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1731.packet_count,1731);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1732.packet_count,1732);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1733.packet_count,1733);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1734.packet_count,1734);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1735.packet_count,1735);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1736.packet_count,1736);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1737.packet_count,1737);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1738.packet_count,1738);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1739.packet_count,1739);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1740.packet_count,1740);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1741.packet_count,1741);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1742.packet_count,1742);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1743.packet_count,1743);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1744.packet_count,1744);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1745.packet_count,1745);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1746.packet_count,1746);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1747.packet_count,1747);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1748.packet_count,1748);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1749.packet_count,1749);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1750.packet_count,1750);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1751.packet_count,1751);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1752.packet_count,1752);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1753.packet_count,1753);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1754.packet_count,1754);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1755.packet_count,1755);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1756.packet_count,1756);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1757.packet_count,1757);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1758.packet_count,1758);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1759.packet_count,1759);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1760.packet_count,1760);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1761.packet_count,1761);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1762.packet_count,1762);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1763.packet_count,1763);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1764.packet_count,1764);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1765.packet_count,1765);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1766.packet_count,1766);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1767.packet_count,1767);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1768.packet_count,1768);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1769.packet_count,1769);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1770.packet_count,1770);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1771.packet_count,1771);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1772.packet_count,1772);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1773.packet_count,1773);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1774.packet_count,1774);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1775.packet_count,1775);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1776.packet_count,1776);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1777.packet_count,1777);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1778.packet_count,1778);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1779.packet_count,1779);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1780.packet_count,1780);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1781.packet_count,1781);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1782.packet_count,1782);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1783.packet_count,1783);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1784.packet_count,1784);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1785.packet_count,1785);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1786.packet_count,1786);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1787.packet_count,1787);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1788.packet_count,1788);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1789.packet_count,1789);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1790.packet_count,1790);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1791.packet_count,1791);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1792.packet_count,1792);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1793.packet_count,1793);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1794.packet_count,1794);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1795.packet_count,1795);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1796.packet_count,1796);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1797.packet_count,1797);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1798.packet_count,1798);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1799.packet_count,1799);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1800.packet_count,1800);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1801.packet_count,1801);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1802.packet_count,1802);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1803.packet_count,1803);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1804.packet_count,1804);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1805.packet_count,1805);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1806.packet_count,1806);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1807.packet_count,1807);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1808.packet_count,1808);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1809.packet_count,1809);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1810.packet_count,1810);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1811.packet_count,1811);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1812.packet_count,1812);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1813.packet_count,1813);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1814.packet_count,1814);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1815.packet_count,1815);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1816.packet_count,1816);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1817.packet_count,1817);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1818.packet_count,1818);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1819.packet_count,1819);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1820.packet_count,1820);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1821.packet_count,1821);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1822.packet_count,1822);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1823.packet_count,1823);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1824.packet_count,1824);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1825.packet_count,1825);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1826.packet_count,1826);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1827.packet_count,1827);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1828.packet_count,1828);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1829.packet_count,1829);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1830.packet_count,1830);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1831.packet_count,1831);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1832.packet_count,1832);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1833.packet_count,1833);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1834.packet_count,1834);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1835.packet_count,1835);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1836.packet_count,1836);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1837.packet_count,1837);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1838.packet_count,1838);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1839.packet_count,1839);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1840.packet_count,1840);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1841.packet_count,1841);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1842.packet_count,1842);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1843.packet_count,1843);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1844.packet_count,1844);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1845.packet_count,1845);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1846.packet_count,1846);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1847.packet_count,1847);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1848.packet_count,1848);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1849.packet_count,1849);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1850.packet_count,1850);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1851.packet_count,1851);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1852.packet_count,1852);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1853.packet_count,1853);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1854.packet_count,1854);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1855.packet_count,1855);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1856.packet_count,1856);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1857.packet_count,1857);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1858.packet_count,1858);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1859.packet_count,1859);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1860.packet_count,1860);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1861.packet_count,1861);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1862.packet_count,1862);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1863.packet_count,1863);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1864.packet_count,1864);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1865.packet_count,1865);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1866.packet_count,1866);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1867.packet_count,1867);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1868.packet_count,1868);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1869.packet_count,1869);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1870.packet_count,1870);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1871.packet_count,1871);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1872.packet_count,1872);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1873.packet_count,1873);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1874.packet_count,1874);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1875.packet_count,1875);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1876.packet_count,1876);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1877.packet_count,1877);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1878.packet_count,1878);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1879.packet_count,1879);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1880.packet_count,1880);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1881.packet_count,1881);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1882.packet_count,1882);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1883.packet_count,1883);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1884.packet_count,1884);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1885.packet_count,1885);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1886.packet_count,1886);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1887.packet_count,1887);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1888.packet_count,1888);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1889.packet_count,1889);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1890.packet_count,1890);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1891.packet_count,1891);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1892.packet_count,1892);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1893.packet_count,1893);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1894.packet_count,1894);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1895.packet_count,1895);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1896.packet_count,1896);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1897.packet_count,1897);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1898.packet_count,1898);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1899.packet_count,1899);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1900.packet_count,1900);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1901.packet_count,1901);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1902.packet_count,1902);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1903.packet_count,1903);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1904.packet_count,1904);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1905.packet_count,1905);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1906.packet_count,1906);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1907.packet_count,1907);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1908.packet_count,1908);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1909.packet_count,1909);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1910.packet_count,1910);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1911.packet_count,1911);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1912.packet_count,1912);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1913.packet_count,1913);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1914.packet_count,1914);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1915.packet_count,1915);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1916.packet_count,1916);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1917.packet_count,1917);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1918.packet_count,1918);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1919.packet_count,1919);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1920.packet_count,1920);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1921.packet_count,1921);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1922.packet_count,1922);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1923.packet_count,1923);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1924.packet_count,1924);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1925.packet_count,1925);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1926.packet_count,1926);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1927.packet_count,1927);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1928.packet_count,1928);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1929.packet_count,1929);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1930.packet_count,1930);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1931.packet_count,1931);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1932.packet_count,1932);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1933.packet_count,1933);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1934.packet_count,1934);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1935.packet_count,1935);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1936.packet_count,1936);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1937.packet_count,1937);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1938.packet_count,1938);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1939.packet_count,1939);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1940.packet_count,1940);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1941.packet_count,1941);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1942.packet_count,1942);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1943.packet_count,1943);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1944.packet_count,1944);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1945.packet_count,1945);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1946.packet_count,1946);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1947.packet_count,1947);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1948.packet_count,1948);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1949.packet_count,1949);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1950.packet_count,1950);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1951.packet_count,1951);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1952.packet_count,1952);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1953.packet_count,1953);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1954.packet_count,1954);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1955.packet_count,1955);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1956.packet_count,1956);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1957.packet_count,1957);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1958.packet_count,1958);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1959.packet_count,1959);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1960.packet_count,1960);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1961.packet_count,1961);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1962.packet_count,1962);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1963.packet_count,1963);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1964.packet_count,1964);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1965.packet_count,1965);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1966.packet_count,1966);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1967.packet_count,1967);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1968.packet_count,1968);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1969.packet_count,1969);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1970.packet_count,1970);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1971.packet_count,1971);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1972.packet_count,1972);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1973.packet_count,1973);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1974.packet_count,1974);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1975.packet_count,1975);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1976.packet_count,1976);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1977.packet_count,1977);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1978.packet_count,1978);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1979.packet_count,1979);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1980.packet_count,1980);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1981.packet_count,1981);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1982.packet_count,1982);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1983.packet_count,1983);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1984.packet_count,1984);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1985.packet_count,1985);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1986.packet_count,1986);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1987.packet_count,1987);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1988.packet_count,1988);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1989.packet_count,1989);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1990.packet_count,1990);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1991.packet_count,1991);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1992.packet_count,1992);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1993.packet_count,1993);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1994.packet_count,1994);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1995.packet_count,1995);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1996.packet_count,1996);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1997.packet_count,1997);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1998.packet_count,1998);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_1999.packet_count,1999);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2000.packet_count,2000);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2001.packet_count,2001);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2002.packet_count,2002);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2003.packet_count,2003);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2004.packet_count,2004);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2005.packet_count,2005);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2006.packet_count,2006);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2007.packet_count,2007);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2008.packet_count,2008);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2009.packet_count,2009);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2010.packet_count,2010);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2011.packet_count,2011);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2012.packet_count,2012);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2013.packet_count,2013);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2014.packet_count,2014);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2015.packet_count,2015);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2016.packet_count,2016);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2017.packet_count,2017);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2018.packet_count,2018);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2019.packet_count,2019);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2020.packet_count,2020);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2021.packet_count,2021);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2022.packet_count,2022);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2023.packet_count,2023);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2024.packet_count,2024);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2025.packet_count,2025);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2026.packet_count,2026);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2027.packet_count,2027);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2028.packet_count,2028);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2029.packet_count,2029);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2030.packet_count,2030);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2031.packet_count,2031);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2032.packet_count,2032);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2033.packet_count,2033);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2034.packet_count,2034);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2035.packet_count,2035);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2036.packet_count,2036);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2037.packet_count,2037);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2038.packet_count,2038);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2039.packet_count,2039);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2040.packet_count,2040);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2041.packet_count,2041);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2042.packet_count,2042);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2043.packet_count,2043);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2044.packet_count,2044);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2045.packet_count,2045);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2046.packet_count,2046);
        packet_count_check(packet_count,env.pf_vf_mux_scbd_2047.packet_count,2047);
      `endif  
  endfunction

  function upstream_final_packet_count_check();
      uvm_config_db#(int)::get(null, "", "no_of_trans", packet_count);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_0_up.packet_count,0);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1_up.packet_count,1);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2_up.packet_count,2);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_3_up.packet_count,3);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_4_up.packet_count,4);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_5_up.packet_count,5);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_6_up.packet_count,6);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_7_up.packet_count,7);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_8_up.packet_count,8);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_9_up.packet_count,9);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_10_up.packet_count,10);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_11_up.packet_count,11);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_12_up.packet_count,12);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_13_up.packet_count,13);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_14_up.packet_count,14);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_15_up.packet_count,15);
      `ifdef TB_CONFIG_2
      packet_count_check(packet_count,env.pf_vf_mux_scbd_16_up.packet_count,16);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_17_up.packet_count,17);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_18_up.packet_count,18);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_19_up.packet_count,19);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_20_up.packet_count,20);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_21_up.packet_count,21);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_22_up.packet_count,22);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_23_up.packet_count,23);
      `elsif TB_CONFIG_3
      packet_count_check(packet_count,env.pf_vf_mux_scbd_16_up.packet_count,16);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_17_up.packet_count,17);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_18_up.packet_count,18);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_19_up.packet_count,19);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_20_up.packet_count,20);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_21_up.packet_count,21);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_22_up.packet_count,22);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_23_up.packet_count,23);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_24_up.packet_count,24);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_25_up.packet_count,25);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_26_up.packet_count,26);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_27_up.packet_count,27);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_28_up.packet_count,28);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_29_up.packet_count,29);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_30_up.packet_count,30);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_31_up.packet_count,31);
      `elsif TB_CONFIG_4
      packet_count_check(packet_count,env.pf_vf_mux_scbd_16_up.packet_count,16);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_17_up.packet_count,17);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_18_up.packet_count,18);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_19_up.packet_count,19);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_20_up.packet_count,20);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_21_up.packet_count,21);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_22_up.packet_count,22);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_23_up.packet_count,23);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_24_up.packet_count,24);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_25_up.packet_count,25);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_26_up.packet_count,26);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_27_up.packet_count,27);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_28_up.packet_count,28);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_29_up.packet_count,29);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_30_up.packet_count,30);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_31_up.packet_count,31);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_32_up.packet_count,32);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_33_up.packet_count,33);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_34_up.packet_count,34);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_35_up.packet_count,35);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_36_up.packet_count,36);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_37_up.packet_count,37);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_38_up.packet_count,38);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_39_up.packet_count,39);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_40_up.packet_count,40);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_41_up.packet_count,41);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_42_up.packet_count,42);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_43_up.packet_count,43);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_44_up.packet_count,44);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_45_up.packet_count,45);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_46_up.packet_count,46);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_47_up.packet_count,47);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_48_up.packet_count,48);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_49_up.packet_count,49);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_50_up.packet_count,50);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_51_up.packet_count,51);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_52_up.packet_count,52);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_53_up.packet_count,53);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_54_up.packet_count,54);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_55_up.packet_count,55);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_56_up.packet_count,56);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_57_up.packet_count,57);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_58_up.packet_count,58);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_59_up.packet_count,59);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_60_up.packet_count,60);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_61_up.packet_count,61);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_62_up.packet_count,62);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_63_up.packet_count,63);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_64_up.packet_count,64);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_65_up.packet_count,65);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_66_up.packet_count,66);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_67_up.packet_count,67);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_68_up.packet_count,68);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_69_up.packet_count,69);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_70_up.packet_count,70);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_71_up.packet_count,71);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_72_up.packet_count,72);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_73_up.packet_count,73);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_74_up.packet_count,74);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_75_up.packet_count,75);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_76_up.packet_count,76);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_77_up.packet_count,77);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_78_up.packet_count,78);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_79_up.packet_count,79);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_80_up.packet_count,80);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_81_up.packet_count,81);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_82_up.packet_count,82);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_83_up.packet_count,83);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_84_up.packet_count,84);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_85_up.packet_count,85);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_86_up.packet_count,86);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_87_up.packet_count,87);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_88_up.packet_count,88);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_89_up.packet_count,89);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_90_up.packet_count,90);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_91_up.packet_count,91);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_92_up.packet_count,92);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_93_up.packet_count,93);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_94_up.packet_count,94);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_95_up.packet_count,95);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_96_up.packet_count,96);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_97_up.packet_count,97);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_98_up.packet_count,98);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_99_up.packet_count,99);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_100_up.packet_count,100);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_101_up.packet_count,101);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_102_up.packet_count,102);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_103_up.packet_count,103);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_104_up.packet_count,104);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_105_up.packet_count,105);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_106_up.packet_count,106);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_107_up.packet_count,107);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_108_up.packet_count,108);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_109_up.packet_count,109);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_110_up.packet_count,110);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_111_up.packet_count,111);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_112_up.packet_count,112);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_113_up.packet_count,113);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_114_up.packet_count,114);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_115_up.packet_count,115);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_116_up.packet_count,116);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_117_up.packet_count,117);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_118_up.packet_count,118);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_119_up.packet_count,119);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_120_up.packet_count,120);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_121_up.packet_count,121);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_122_up.packet_count,122);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_123_up.packet_count,123);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_124_up.packet_count,124);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_125_up.packet_count,125);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_126_up.packet_count,126);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_127_up.packet_count,127);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_128_up.packet_count,128);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_129_up.packet_count,129);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_130_up.packet_count,130);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_131_up.packet_count,131);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_132_up.packet_count,132);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_133_up.packet_count,133);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_134_up.packet_count,134);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_135_up.packet_count,135);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_136_up.packet_count,136);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_137_up.packet_count,137);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_138_up.packet_count,138);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_139_up.packet_count,139);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_140_up.packet_count,140);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_141_up.packet_count,141);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_142_up.packet_count,142);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_143_up.packet_count,143);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_144_up.packet_count,144);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_145_up.packet_count,145);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_146_up.packet_count,146);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_147_up.packet_count,147);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_148_up.packet_count,148);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_149_up.packet_count,149);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_150_up.packet_count,150);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_151_up.packet_count,151);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_152_up.packet_count,152);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_153_up.packet_count,153);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_154_up.packet_count,154);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_155_up.packet_count,155);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_156_up.packet_count,156);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_157_up.packet_count,157);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_158_up.packet_count,158);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_159_up.packet_count,159);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_160_up.packet_count,160);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_161_up.packet_count,161);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_162_up.packet_count,162);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_163_up.packet_count,163);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_164_up.packet_count,164);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_165_up.packet_count,165);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_166_up.packet_count,166);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_167_up.packet_count,167);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_168_up.packet_count,168);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_169_up.packet_count,169);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_170_up.packet_count,170);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_171_up.packet_count,171);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_172_up.packet_count,172);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_173_up.packet_count,173);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_174_up.packet_count,174);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_175_up.packet_count,175);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_176_up.packet_count,176);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_177_up.packet_count,177);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_178_up.packet_count,178);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_179_up.packet_count,179);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_180_up.packet_count,180);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_181_up.packet_count,181);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_182_up.packet_count,182);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_183_up.packet_count,183);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_184_up.packet_count,184);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_185_up.packet_count,185);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_186_up.packet_count,186);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_187_up.packet_count,187);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_188_up.packet_count,188);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_189_up.packet_count,189);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_190_up.packet_count,190);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_191_up.packet_count,191);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_192_up.packet_count,192);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_193_up.packet_count,193);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_194_up.packet_count,194);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_195_up.packet_count,195);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_196_up.packet_count,196);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_197_up.packet_count,197);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_198_up.packet_count,198);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_199_up.packet_count,199);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_200_up.packet_count,200);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_201_up.packet_count,201);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_202_up.packet_count,202);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_203_up.packet_count,203);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_204_up.packet_count,204);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_205_up.packet_count,205);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_206_up.packet_count,206);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_207_up.packet_count,207);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_208_up.packet_count,208);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_209_up.packet_count,209);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_210_up.packet_count,210);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_211_up.packet_count,211);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_212_up.packet_count,212);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_213_up.packet_count,213);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_214_up.packet_count,214);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_215_up.packet_count,215);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_216_up.packet_count,216);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_217_up.packet_count,217);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_218_up.packet_count,218);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_219_up.packet_count,219);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_220_up.packet_count,220);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_221_up.packet_count,221);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_222_up.packet_count,222);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_223_up.packet_count,223);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_224_up.packet_count,224);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_225_up.packet_count,225);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_226_up.packet_count,226);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_227_up.packet_count,227);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_228_up.packet_count,228);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_229_up.packet_count,229);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_230_up.packet_count,230);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_231_up.packet_count,231);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_232_up.packet_count,232);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_233_up.packet_count,233);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_234_up.packet_count,234);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_235_up.packet_count,235);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_236_up.packet_count,236);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_237_up.packet_count,237);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_238_up.packet_count,238);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_239_up.packet_count,239);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_240_up.packet_count,240);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_241_up.packet_count,241);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_242_up.packet_count,242);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_243_up.packet_count,243);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_244_up.packet_count,244);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_245_up.packet_count,245);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_246_up.packet_count,246);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_247_up.packet_count,247);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_248_up.packet_count,248);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_249_up.packet_count,249);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_250_up.packet_count,250);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_251_up.packet_count,251);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_252_up.packet_count,252);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_253_up.packet_count,253);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_254_up.packet_count,254);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_255_up.packet_count,255);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_256_up.packet_count,256);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_257_up.packet_count,257);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_258_up.packet_count,258);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_259_up.packet_count,259);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_260_up.packet_count,260);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_261_up.packet_count,261);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_262_up.packet_count,262);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_263_up.packet_count,263);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_264_up.packet_count,264);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_265_up.packet_count,265);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_266_up.packet_count,266);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_267_up.packet_count,267);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_268_up.packet_count,268);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_269_up.packet_count,269);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_270_up.packet_count,270);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_271_up.packet_count,271);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_272_up.packet_count,272);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_273_up.packet_count,273);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_274_up.packet_count,274);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_275_up.packet_count,275);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_276_up.packet_count,276);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_277_up.packet_count,277);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_278_up.packet_count,278);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_279_up.packet_count,279);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_280_up.packet_count,280);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_281_up.packet_count,281);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_282_up.packet_count,282);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_283_up.packet_count,283);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_284_up.packet_count,284);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_285_up.packet_count,285);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_286_up.packet_count,286);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_287_up.packet_count,287);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_288_up.packet_count,288);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_289_up.packet_count,289);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_290_up.packet_count,290);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_291_up.packet_count,291);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_292_up.packet_count,292);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_293_up.packet_count,293);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_294_up.packet_count,294);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_295_up.packet_count,295);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_296_up.packet_count,296);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_297_up.packet_count,297);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_298_up.packet_count,298);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_299_up.packet_count,299);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_300_up.packet_count,300);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_301_up.packet_count,301);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_302_up.packet_count,302);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_303_up.packet_count,303);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_304_up.packet_count,304);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_305_up.packet_count,305);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_306_up.packet_count,306);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_307_up.packet_count,307);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_308_up.packet_count,308);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_309_up.packet_count,309);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_310_up.packet_count,310);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_311_up.packet_count,311);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_312_up.packet_count,312);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_313_up.packet_count,313);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_314_up.packet_count,314);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_315_up.packet_count,315);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_316_up.packet_count,316);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_317_up.packet_count,317);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_318_up.packet_count,318);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_319_up.packet_count,319);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_320_up.packet_count,320);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_321_up.packet_count,321);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_322_up.packet_count,322);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_323_up.packet_count,323);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_324_up.packet_count,324);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_325_up.packet_count,325);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_326_up.packet_count,326);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_327_up.packet_count,327);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_328_up.packet_count,328);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_329_up.packet_count,329);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_330_up.packet_count,330);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_331_up.packet_count,331);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_332_up.packet_count,332);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_333_up.packet_count,333);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_334_up.packet_count,334);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_335_up.packet_count,335);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_336_up.packet_count,336);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_337_up.packet_count,337);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_338_up.packet_count,338);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_339_up.packet_count,339);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_340_up.packet_count,340);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_341_up.packet_count,341);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_342_up.packet_count,342);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_343_up.packet_count,343);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_344_up.packet_count,344);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_345_up.packet_count,345);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_346_up.packet_count,346);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_347_up.packet_count,347);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_348_up.packet_count,348);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_349_up.packet_count,349);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_350_up.packet_count,350);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_351_up.packet_count,351);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_352_up.packet_count,352);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_353_up.packet_count,353);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_354_up.packet_count,354);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_355_up.packet_count,355);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_356_up.packet_count,356);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_357_up.packet_count,357);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_358_up.packet_count,358);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_359_up.packet_count,359);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_360_up.packet_count,360);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_361_up.packet_count,361);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_362_up.packet_count,362);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_363_up.packet_count,363);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_364_up.packet_count,364);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_365_up.packet_count,365);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_366_up.packet_count,366);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_367_up.packet_count,367);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_368_up.packet_count,368);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_369_up.packet_count,369);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_370_up.packet_count,370);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_371_up.packet_count,371);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_372_up.packet_count,372);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_373_up.packet_count,373);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_374_up.packet_count,374);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_375_up.packet_count,375);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_376_up.packet_count,376);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_377_up.packet_count,377);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_378_up.packet_count,378);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_379_up.packet_count,379);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_380_up.packet_count,380);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_381_up.packet_count,381);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_382_up.packet_count,382);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_383_up.packet_count,383);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_384_up.packet_count,384);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_385_up.packet_count,385);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_386_up.packet_count,386);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_387_up.packet_count,387);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_388_up.packet_count,388);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_389_up.packet_count,389);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_390_up.packet_count,390);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_391_up.packet_count,391);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_392_up.packet_count,392);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_393_up.packet_count,393);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_394_up.packet_count,394);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_395_up.packet_count,395);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_396_up.packet_count,396);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_397_up.packet_count,397);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_398_up.packet_count,398);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_399_up.packet_count,399);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_400_up.packet_count,400);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_401_up.packet_count,401);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_402_up.packet_count,402);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_403_up.packet_count,403);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_404_up.packet_count,404);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_405_up.packet_count,405);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_406_up.packet_count,406);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_407_up.packet_count,407);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_408_up.packet_count,408);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_409_up.packet_count,409);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_410_up.packet_count,410);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_411_up.packet_count,411);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_412_up.packet_count,412);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_413_up.packet_count,413);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_414_up.packet_count,414);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_415_up.packet_count,415);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_416_up.packet_count,416);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_417_up.packet_count,417);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_418_up.packet_count,418);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_419_up.packet_count,419);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_420_up.packet_count,420);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_421_up.packet_count,421);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_422_up.packet_count,422);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_423_up.packet_count,423);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_424_up.packet_count,424);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_425_up.packet_count,425);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_426_up.packet_count,426);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_427_up.packet_count,427);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_428_up.packet_count,428);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_429_up.packet_count,429);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_430_up.packet_count,430);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_431_up.packet_count,431);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_432_up.packet_count,432);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_433_up.packet_count,433);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_434_up.packet_count,434);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_435_up.packet_count,435);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_436_up.packet_count,436);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_437_up.packet_count,437);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_438_up.packet_count,438);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_439_up.packet_count,439);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_440_up.packet_count,440);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_441_up.packet_count,441);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_442_up.packet_count,442);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_443_up.packet_count,443);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_444_up.packet_count,444);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_445_up.packet_count,445);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_446_up.packet_count,446);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_447_up.packet_count,447);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_448_up.packet_count,448);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_449_up.packet_count,449);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_450_up.packet_count,450);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_451_up.packet_count,451);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_452_up.packet_count,452);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_453_up.packet_count,453);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_454_up.packet_count,454);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_455_up.packet_count,455);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_456_up.packet_count,456);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_457_up.packet_count,457);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_458_up.packet_count,458);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_459_up.packet_count,459);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_460_up.packet_count,460);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_461_up.packet_count,461);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_462_up.packet_count,462);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_463_up.packet_count,463);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_464_up.packet_count,464);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_465_up.packet_count,465);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_466_up.packet_count,466);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_467_up.packet_count,467);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_468_up.packet_count,468);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_469_up.packet_count,469);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_470_up.packet_count,470);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_471_up.packet_count,471);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_472_up.packet_count,472);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_473_up.packet_count,473);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_474_up.packet_count,474);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_475_up.packet_count,475);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_476_up.packet_count,476);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_477_up.packet_count,477);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_478_up.packet_count,478);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_479_up.packet_count,479);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_480_up.packet_count,480);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_481_up.packet_count,481);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_482_up.packet_count,482);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_483_up.packet_count,483);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_484_up.packet_count,484);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_485_up.packet_count,485);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_486_up.packet_count,486);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_487_up.packet_count,487);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_488_up.packet_count,488);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_489_up.packet_count,489);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_490_up.packet_count,490);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_491_up.packet_count,491);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_492_up.packet_count,492);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_493_up.packet_count,493);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_494_up.packet_count,494);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_495_up.packet_count,495);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_496_up.packet_count,496);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_497_up.packet_count,497);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_498_up.packet_count,498);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_499_up.packet_count,499);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_500_up.packet_count,500);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_501_up.packet_count,501);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_502_up.packet_count,502);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_503_up.packet_count,503);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_504_up.packet_count,504);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_505_up.packet_count,505);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_506_up.packet_count,506);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_507_up.packet_count,507);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_508_up.packet_count,508);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_509_up.packet_count,509);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_510_up.packet_count,510);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_511_up.packet_count,511);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_512_up.packet_count,512);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_513_up.packet_count,513);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_514_up.packet_count,514);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_515_up.packet_count,515);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_516_up.packet_count,516);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_517_up.packet_count,517);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_518_up.packet_count,518);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_519_up.packet_count,519);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_520_up.packet_count,520);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_521_up.packet_count,521);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_522_up.packet_count,522);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_523_up.packet_count,523);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_524_up.packet_count,524);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_525_up.packet_count,525);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_526_up.packet_count,526);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_527_up.packet_count,527);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_528_up.packet_count,528);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_529_up.packet_count,529);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_530_up.packet_count,530);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_531_up.packet_count,531);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_532_up.packet_count,532);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_533_up.packet_count,533);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_534_up.packet_count,534);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_535_up.packet_count,535);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_536_up.packet_count,536);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_537_up.packet_count,537);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_538_up.packet_count,538);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_539_up.packet_count,539);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_540_up.packet_count,540);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_541_up.packet_count,541);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_542_up.packet_count,542);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_543_up.packet_count,543);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_544_up.packet_count,544);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_545_up.packet_count,545);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_546_up.packet_count,546);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_547_up.packet_count,547);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_548_up.packet_count,548);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_549_up.packet_count,549);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_550_up.packet_count,550);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_551_up.packet_count,551);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_552_up.packet_count,552);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_553_up.packet_count,553);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_554_up.packet_count,554);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_555_up.packet_count,555);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_556_up.packet_count,556);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_557_up.packet_count,557);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_558_up.packet_count,558);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_559_up.packet_count,559);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_560_up.packet_count,560);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_561_up.packet_count,561);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_562_up.packet_count,562);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_563_up.packet_count,563);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_564_up.packet_count,564);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_565_up.packet_count,565);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_566_up.packet_count,566);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_567_up.packet_count,567);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_568_up.packet_count,568);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_569_up.packet_count,569);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_570_up.packet_count,570);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_571_up.packet_count,571);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_572_up.packet_count,572);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_573_up.packet_count,573);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_574_up.packet_count,574);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_575_up.packet_count,575);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_576_up.packet_count,576);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_577_up.packet_count,577);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_578_up.packet_count,578);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_579_up.packet_count,579);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_580_up.packet_count,580);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_581_up.packet_count,581);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_582_up.packet_count,582);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_583_up.packet_count,583);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_584_up.packet_count,584);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_585_up.packet_count,585);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_586_up.packet_count,586);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_587_up.packet_count,587);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_588_up.packet_count,588);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_589_up.packet_count,589);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_590_up.packet_count,590);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_591_up.packet_count,591);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_592_up.packet_count,592);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_593_up.packet_count,593);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_594_up.packet_count,594);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_595_up.packet_count,595);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_596_up.packet_count,596);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_597_up.packet_count,597);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_598_up.packet_count,598);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_599_up.packet_count,599);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_600_up.packet_count,600);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_601_up.packet_count,601);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_602_up.packet_count,602);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_603_up.packet_count,603);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_604_up.packet_count,604);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_605_up.packet_count,605);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_606_up.packet_count,606);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_607_up.packet_count,607);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_608_up.packet_count,608);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_609_up.packet_count,609);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_610_up.packet_count,610);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_611_up.packet_count,611);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_612_up.packet_count,612);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_613_up.packet_count,613);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_614_up.packet_count,614);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_615_up.packet_count,615);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_616_up.packet_count,616);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_617_up.packet_count,617);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_618_up.packet_count,618);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_619_up.packet_count,619);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_620_up.packet_count,620);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_621_up.packet_count,621);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_622_up.packet_count,622);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_623_up.packet_count,623);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_624_up.packet_count,624);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_625_up.packet_count,625);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_626_up.packet_count,626);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_627_up.packet_count,627);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_628_up.packet_count,628);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_629_up.packet_count,629);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_630_up.packet_count,630);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_631_up.packet_count,631);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_632_up.packet_count,632);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_633_up.packet_count,633);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_634_up.packet_count,634);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_635_up.packet_count,635);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_636_up.packet_count,636);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_637_up.packet_count,637);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_638_up.packet_count,638);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_639_up.packet_count,639);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_640_up.packet_count,640);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_641_up.packet_count,641);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_642_up.packet_count,642);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_643_up.packet_count,643);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_644_up.packet_count,644);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_645_up.packet_count,645);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_646_up.packet_count,646);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_647_up.packet_count,647);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_648_up.packet_count,648);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_649_up.packet_count,649);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_650_up.packet_count,650);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_651_up.packet_count,651);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_652_up.packet_count,652);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_653_up.packet_count,653);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_654_up.packet_count,654);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_655_up.packet_count,655);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_656_up.packet_count,656);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_657_up.packet_count,657);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_658_up.packet_count,658);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_659_up.packet_count,659);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_660_up.packet_count,660);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_661_up.packet_count,661);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_662_up.packet_count,662);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_663_up.packet_count,663);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_664_up.packet_count,664);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_665_up.packet_count,665);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_666_up.packet_count,666);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_667_up.packet_count,667);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_668_up.packet_count,668);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_669_up.packet_count,669);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_670_up.packet_count,670);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_671_up.packet_count,671);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_672_up.packet_count,672);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_673_up.packet_count,673);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_674_up.packet_count,674);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_675_up.packet_count,675);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_676_up.packet_count,676);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_677_up.packet_count,677);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_678_up.packet_count,678);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_679_up.packet_count,679);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_680_up.packet_count,680);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_681_up.packet_count,681);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_682_up.packet_count,682);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_683_up.packet_count,683);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_684_up.packet_count,684);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_685_up.packet_count,685);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_686_up.packet_count,686);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_687_up.packet_count,687);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_688_up.packet_count,688);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_689_up.packet_count,689);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_690_up.packet_count,690);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_691_up.packet_count,691);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_692_up.packet_count,692);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_693_up.packet_count,693);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_694_up.packet_count,694);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_695_up.packet_count,695);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_696_up.packet_count,696);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_697_up.packet_count,697);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_698_up.packet_count,698);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_699_up.packet_count,699);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_700_up.packet_count,700);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_701_up.packet_count,701);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_702_up.packet_count,702);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_703_up.packet_count,703);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_704_up.packet_count,704);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_705_up.packet_count,705);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_706_up.packet_count,706);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_707_up.packet_count,707);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_708_up.packet_count,708);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_709_up.packet_count,709);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_710_up.packet_count,710);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_711_up.packet_count,711);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_712_up.packet_count,712);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_713_up.packet_count,713);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_714_up.packet_count,714);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_715_up.packet_count,715);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_716_up.packet_count,716);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_717_up.packet_count,717);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_718_up.packet_count,718);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_719_up.packet_count,719);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_720_up.packet_count,720);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_721_up.packet_count,721);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_722_up.packet_count,722);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_723_up.packet_count,723);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_724_up.packet_count,724);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_725_up.packet_count,725);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_726_up.packet_count,726);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_727_up.packet_count,727);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_728_up.packet_count,728);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_729_up.packet_count,729);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_730_up.packet_count,730);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_731_up.packet_count,731);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_732_up.packet_count,732);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_733_up.packet_count,733);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_734_up.packet_count,734);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_735_up.packet_count,735);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_736_up.packet_count,736);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_737_up.packet_count,737);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_738_up.packet_count,738);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_739_up.packet_count,739);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_740_up.packet_count,740);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_741_up.packet_count,741);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_742_up.packet_count,742);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_743_up.packet_count,743);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_744_up.packet_count,744);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_745_up.packet_count,745);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_746_up.packet_count,746);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_747_up.packet_count,747);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_748_up.packet_count,748);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_749_up.packet_count,749);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_750_up.packet_count,750);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_751_up.packet_count,751);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_752_up.packet_count,752);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_753_up.packet_count,753);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_754_up.packet_count,754);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_755_up.packet_count,755);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_756_up.packet_count,756);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_757_up.packet_count,757);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_758_up.packet_count,758);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_759_up.packet_count,759);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_760_up.packet_count,760);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_761_up.packet_count,761);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_762_up.packet_count,762);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_763_up.packet_count,763);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_764_up.packet_count,764);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_765_up.packet_count,765);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_766_up.packet_count,766);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_767_up.packet_count,767);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_768_up.packet_count,768);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_769_up.packet_count,769);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_770_up.packet_count,770);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_771_up.packet_count,771);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_772_up.packet_count,772);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_773_up.packet_count,773);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_774_up.packet_count,774);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_775_up.packet_count,775);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_776_up.packet_count,776);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_777_up.packet_count,777);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_778_up.packet_count,778);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_779_up.packet_count,779);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_780_up.packet_count,780);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_781_up.packet_count,781);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_782_up.packet_count,782);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_783_up.packet_count,783);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_784_up.packet_count,784);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_785_up.packet_count,785);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_786_up.packet_count,786);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_787_up.packet_count,787);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_788_up.packet_count,788);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_789_up.packet_count,789);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_790_up.packet_count,790);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_791_up.packet_count,791);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_792_up.packet_count,792);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_793_up.packet_count,793);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_794_up.packet_count,794);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_795_up.packet_count,795);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_796_up.packet_count,796);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_797_up.packet_count,797);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_798_up.packet_count,798);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_799_up.packet_count,799);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_800_up.packet_count,800);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_801_up.packet_count,801);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_802_up.packet_count,802);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_803_up.packet_count,803);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_804_up.packet_count,804);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_805_up.packet_count,805);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_806_up.packet_count,806);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_807_up.packet_count,807);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_808_up.packet_count,808);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_809_up.packet_count,809);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_810_up.packet_count,810);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_811_up.packet_count,811);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_812_up.packet_count,812);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_813_up.packet_count,813);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_814_up.packet_count,814);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_815_up.packet_count,815);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_816_up.packet_count,816);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_817_up.packet_count,817);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_818_up.packet_count,818);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_819_up.packet_count,819);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_820_up.packet_count,820);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_821_up.packet_count,821);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_822_up.packet_count,822);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_823_up.packet_count,823);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_824_up.packet_count,824);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_825_up.packet_count,825);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_826_up.packet_count,826);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_827_up.packet_count,827);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_828_up.packet_count,828);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_829_up.packet_count,829);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_830_up.packet_count,830);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_831_up.packet_count,831);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_832_up.packet_count,832);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_833_up.packet_count,833);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_834_up.packet_count,834);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_835_up.packet_count,835);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_836_up.packet_count,836);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_837_up.packet_count,837);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_838_up.packet_count,838);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_839_up.packet_count,839);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_840_up.packet_count,840);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_841_up.packet_count,841);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_842_up.packet_count,842);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_843_up.packet_count,843);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_844_up.packet_count,844);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_845_up.packet_count,845);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_846_up.packet_count,846);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_847_up.packet_count,847);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_848_up.packet_count,848);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_849_up.packet_count,849);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_850_up.packet_count,850);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_851_up.packet_count,851);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_852_up.packet_count,852);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_853_up.packet_count,853);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_854_up.packet_count,854);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_855_up.packet_count,855);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_856_up.packet_count,856);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_857_up.packet_count,857);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_858_up.packet_count,858);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_859_up.packet_count,859);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_860_up.packet_count,860);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_861_up.packet_count,861);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_862_up.packet_count,862);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_863_up.packet_count,863);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_864_up.packet_count,864);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_865_up.packet_count,865);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_866_up.packet_count,866);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_867_up.packet_count,867);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_868_up.packet_count,868);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_869_up.packet_count,869);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_870_up.packet_count,870);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_871_up.packet_count,871);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_872_up.packet_count,872);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_873_up.packet_count,873);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_874_up.packet_count,874);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_875_up.packet_count,875);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_876_up.packet_count,876);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_877_up.packet_count,877);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_878_up.packet_count,878);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_879_up.packet_count,879);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_880_up.packet_count,880);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_881_up.packet_count,881);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_882_up.packet_count,882);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_883_up.packet_count,883);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_884_up.packet_count,884);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_885_up.packet_count,885);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_886_up.packet_count,886);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_887_up.packet_count,887);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_888_up.packet_count,888);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_889_up.packet_count,889);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_890_up.packet_count,890);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_891_up.packet_count,891);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_892_up.packet_count,892);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_893_up.packet_count,893);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_894_up.packet_count,894);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_895_up.packet_count,895);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_896_up.packet_count,896);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_897_up.packet_count,897);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_898_up.packet_count,898);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_899_up.packet_count,899);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_900_up.packet_count,900);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_901_up.packet_count,901);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_902_up.packet_count,902);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_903_up.packet_count,903);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_904_up.packet_count,904);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_905_up.packet_count,905);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_906_up.packet_count,906);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_907_up.packet_count,907);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_908_up.packet_count,908);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_909_up.packet_count,909);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_910_up.packet_count,910);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_911_up.packet_count,911);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_912_up.packet_count,912);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_913_up.packet_count,913);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_914_up.packet_count,914);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_915_up.packet_count,915);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_916_up.packet_count,916);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_917_up.packet_count,917);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_918_up.packet_count,918);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_919_up.packet_count,919);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_920_up.packet_count,920);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_921_up.packet_count,921);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_922_up.packet_count,922);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_923_up.packet_count,923);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_924_up.packet_count,924);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_925_up.packet_count,925);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_926_up.packet_count,926);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_927_up.packet_count,927);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_928_up.packet_count,928);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_929_up.packet_count,929);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_930_up.packet_count,930);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_931_up.packet_count,931);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_932_up.packet_count,932);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_933_up.packet_count,933);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_934_up.packet_count,934);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_935_up.packet_count,935);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_936_up.packet_count,936);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_937_up.packet_count,937);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_938_up.packet_count,938);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_939_up.packet_count,939);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_940_up.packet_count,940);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_941_up.packet_count,941);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_942_up.packet_count,942);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_943_up.packet_count,943);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_944_up.packet_count,944);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_945_up.packet_count,945);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_946_up.packet_count,946);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_947_up.packet_count,947);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_948_up.packet_count,948);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_949_up.packet_count,949);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_950_up.packet_count,950);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_951_up.packet_count,951);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_952_up.packet_count,952);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_953_up.packet_count,953);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_954_up.packet_count,954);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_955_up.packet_count,955);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_956_up.packet_count,956);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_957_up.packet_count,957);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_958_up.packet_count,958);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_959_up.packet_count,959);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_960_up.packet_count,960);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_961_up.packet_count,961);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_962_up.packet_count,962);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_963_up.packet_count,963);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_964_up.packet_count,964);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_965_up.packet_count,965);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_966_up.packet_count,966);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_967_up.packet_count,967);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_968_up.packet_count,968);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_969_up.packet_count,969);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_970_up.packet_count,970);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_971_up.packet_count,971);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_972_up.packet_count,972);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_973_up.packet_count,973);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_974_up.packet_count,974);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_975_up.packet_count,975);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_976_up.packet_count,976);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_977_up.packet_count,977);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_978_up.packet_count,978);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_979_up.packet_count,979);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_980_up.packet_count,980);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_981_up.packet_count,981);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_982_up.packet_count,982);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_983_up.packet_count,983);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_984_up.packet_count,984);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_985_up.packet_count,985);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_986_up.packet_count,986);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_987_up.packet_count,987);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_988_up.packet_count,988);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_989_up.packet_count,989);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_990_up.packet_count,990);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_991_up.packet_count,991);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_992_up.packet_count,992);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_993_up.packet_count,993);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_994_up.packet_count,994);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_995_up.packet_count,995);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_996_up.packet_count,996);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_997_up.packet_count,997);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_998_up.packet_count,998);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_999_up.packet_count,999);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1000_up.packet_count,1000);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1001_up.packet_count,1001);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1002_up.packet_count,1002);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1003_up.packet_count,1003);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1004_up.packet_count,1004);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1005_up.packet_count,1005);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1006_up.packet_count,1006);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1007_up.packet_count,1007);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1008_up.packet_count,1008);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1009_up.packet_count,1009);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1010_up.packet_count,1010);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1011_up.packet_count,1011);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1012_up.packet_count,1012);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1013_up.packet_count,1013);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1014_up.packet_count,1014);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1015_up.packet_count,1015);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1016_up.packet_count,1016);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1017_up.packet_count,1017);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1018_up.packet_count,1018);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1019_up.packet_count,1019);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1020_up.packet_count,1020);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1021_up.packet_count,1021);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1022_up.packet_count,1022);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1023_up.packet_count,1023);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1024_up.packet_count,1024);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1025_up.packet_count,1025);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1026_up.packet_count,1026);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1027_up.packet_count,1027);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1028_up.packet_count,1028);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1029_up.packet_count,1029);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1030_up.packet_count,1030);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1031_up.packet_count,1031);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1032_up.packet_count,1032);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1033_up.packet_count,1033);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1034_up.packet_count,1034);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1035_up.packet_count,1035);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1036_up.packet_count,1036);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1037_up.packet_count,1037);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1038_up.packet_count,1038);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1039_up.packet_count,1039);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1040_up.packet_count,1040);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1041_up.packet_count,1041);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1042_up.packet_count,1042);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1043_up.packet_count,1043);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1044_up.packet_count,1044);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1045_up.packet_count,1045);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1046_up.packet_count,1046);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1047_up.packet_count,1047);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1048_up.packet_count,1048);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1049_up.packet_count,1049);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1050_up.packet_count,1050);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1051_up.packet_count,1051);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1052_up.packet_count,1052);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1053_up.packet_count,1053);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1054_up.packet_count,1054);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1055_up.packet_count,1055);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1056_up.packet_count,1056);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1057_up.packet_count,1057);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1058_up.packet_count,1058);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1059_up.packet_count,1059);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1060_up.packet_count,1060);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1061_up.packet_count,1061);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1062_up.packet_count,1062);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1063_up.packet_count,1063);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1064_up.packet_count,1064);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1065_up.packet_count,1065);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1066_up.packet_count,1066);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1067_up.packet_count,1067);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1068_up.packet_count,1068);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1069_up.packet_count,1069);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1070_up.packet_count,1070);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1071_up.packet_count,1071);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1072_up.packet_count,1072);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1073_up.packet_count,1073);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1074_up.packet_count,1074);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1075_up.packet_count,1075);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1076_up.packet_count,1076);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1077_up.packet_count,1077);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1078_up.packet_count,1078);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1079_up.packet_count,1079);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1080_up.packet_count,1080);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1081_up.packet_count,1081);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1082_up.packet_count,1082);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1083_up.packet_count,1083);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1084_up.packet_count,1084);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1085_up.packet_count,1085);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1086_up.packet_count,1086);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1087_up.packet_count,1087);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1088_up.packet_count,1088);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1089_up.packet_count,1089);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1090_up.packet_count,1090);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1091_up.packet_count,1091);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1092_up.packet_count,1092);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1093_up.packet_count,1093);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1094_up.packet_count,1094);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1095_up.packet_count,1095);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1096_up.packet_count,1096);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1097_up.packet_count,1097);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1098_up.packet_count,1098);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1099_up.packet_count,1099);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1100_up.packet_count,1100);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1101_up.packet_count,1101);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1102_up.packet_count,1102);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1103_up.packet_count,1103);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1104_up.packet_count,1104);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1105_up.packet_count,1105);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1106_up.packet_count,1106);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1107_up.packet_count,1107);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1108_up.packet_count,1108);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1109_up.packet_count,1109);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1110_up.packet_count,1110);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1111_up.packet_count,1111);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1112_up.packet_count,1112);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1113_up.packet_count,1113);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1114_up.packet_count,1114);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1115_up.packet_count,1115);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1116_up.packet_count,1116);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1117_up.packet_count,1117);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1118_up.packet_count,1118);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1119_up.packet_count,1119);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1120_up.packet_count,1120);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1121_up.packet_count,1121);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1122_up.packet_count,1122);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1123_up.packet_count,1123);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1124_up.packet_count,1124);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1125_up.packet_count,1125);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1126_up.packet_count,1126);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1127_up.packet_count,1127);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1128_up.packet_count,1128);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1129_up.packet_count,1129);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1130_up.packet_count,1130);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1131_up.packet_count,1131);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1132_up.packet_count,1132);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1133_up.packet_count,1133);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1134_up.packet_count,1134);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1135_up.packet_count,1135);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1136_up.packet_count,1136);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1137_up.packet_count,1137);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1138_up.packet_count,1138);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1139_up.packet_count,1139);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1140_up.packet_count,1140);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1141_up.packet_count,1141);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1142_up.packet_count,1142);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1143_up.packet_count,1143);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1144_up.packet_count,1144);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1145_up.packet_count,1145);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1146_up.packet_count,1146);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1147_up.packet_count,1147);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1148_up.packet_count,1148);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1149_up.packet_count,1149);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1150_up.packet_count,1150);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1151_up.packet_count,1151);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1152_up.packet_count,1152);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1153_up.packet_count,1153);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1154_up.packet_count,1154);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1155_up.packet_count,1155);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1156_up.packet_count,1156);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1157_up.packet_count,1157);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1158_up.packet_count,1158);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1159_up.packet_count,1159);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1160_up.packet_count,1160);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1161_up.packet_count,1161);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1162_up.packet_count,1162);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1163_up.packet_count,1163);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1164_up.packet_count,1164);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1165_up.packet_count,1165);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1166_up.packet_count,1166);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1167_up.packet_count,1167);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1168_up.packet_count,1168);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1169_up.packet_count,1169);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1170_up.packet_count,1170);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1171_up.packet_count,1171);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1172_up.packet_count,1172);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1173_up.packet_count,1173);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1174_up.packet_count,1174);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1175_up.packet_count,1175);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1176_up.packet_count,1176);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1177_up.packet_count,1177);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1178_up.packet_count,1178);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1179_up.packet_count,1179);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1180_up.packet_count,1180);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1181_up.packet_count,1181);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1182_up.packet_count,1182);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1183_up.packet_count,1183);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1184_up.packet_count,1184);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1185_up.packet_count,1185);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1186_up.packet_count,1186);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1187_up.packet_count,1187);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1188_up.packet_count,1188);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1189_up.packet_count,1189);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1190_up.packet_count,1190);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1191_up.packet_count,1191);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1192_up.packet_count,1192);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1193_up.packet_count,1193);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1194_up.packet_count,1194);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1195_up.packet_count,1195);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1196_up.packet_count,1196);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1197_up.packet_count,1197);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1198_up.packet_count,1198);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1199_up.packet_count,1199);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1200_up.packet_count,1200);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1201_up.packet_count,1201);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1202_up.packet_count,1202);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1203_up.packet_count,1203);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1204_up.packet_count,1204);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1205_up.packet_count,1205);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1206_up.packet_count,1206);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1207_up.packet_count,1207);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1208_up.packet_count,1208);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1209_up.packet_count,1209);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1210_up.packet_count,1210);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1211_up.packet_count,1211);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1212_up.packet_count,1212);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1213_up.packet_count,1213);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1214_up.packet_count,1214);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1215_up.packet_count,1215);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1216_up.packet_count,1216);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1217_up.packet_count,1217);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1218_up.packet_count,1218);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1219_up.packet_count,1219);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1220_up.packet_count,1220);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1221_up.packet_count,1221);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1222_up.packet_count,1222);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1223_up.packet_count,1223);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1224_up.packet_count,1224);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1225_up.packet_count,1225);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1226_up.packet_count,1226);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1227_up.packet_count,1227);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1228_up.packet_count,1228);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1229_up.packet_count,1229);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1230_up.packet_count,1230);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1231_up.packet_count,1231);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1232_up.packet_count,1232);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1233_up.packet_count,1233);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1234_up.packet_count,1234);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1235_up.packet_count,1235);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1236_up.packet_count,1236);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1237_up.packet_count,1237);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1238_up.packet_count,1238);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1239_up.packet_count,1239);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1240_up.packet_count,1240);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1241_up.packet_count,1241);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1242_up.packet_count,1242);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1243_up.packet_count,1243);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1244_up.packet_count,1244);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1245_up.packet_count,1245);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1246_up.packet_count,1246);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1247_up.packet_count,1247);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1248_up.packet_count,1248);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1249_up.packet_count,1249);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1250_up.packet_count,1250);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1251_up.packet_count,1251);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1252_up.packet_count,1252);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1253_up.packet_count,1253);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1254_up.packet_count,1254);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1255_up.packet_count,1255);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1256_up.packet_count,1256);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1257_up.packet_count,1257);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1258_up.packet_count,1258);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1259_up.packet_count,1259);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1260_up.packet_count,1260);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1261_up.packet_count,1261);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1262_up.packet_count,1262);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1263_up.packet_count,1263);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1264_up.packet_count,1264);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1265_up.packet_count,1265);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1266_up.packet_count,1266);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1267_up.packet_count,1267);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1268_up.packet_count,1268);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1269_up.packet_count,1269);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1270_up.packet_count,1270);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1271_up.packet_count,1271);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1272_up.packet_count,1272);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1273_up.packet_count,1273);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1274_up.packet_count,1274);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1275_up.packet_count,1275);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1276_up.packet_count,1276);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1277_up.packet_count,1277);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1278_up.packet_count,1278);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1279_up.packet_count,1279);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1280_up.packet_count,1280);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1281_up.packet_count,1281);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1282_up.packet_count,1282);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1283_up.packet_count,1283);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1284_up.packet_count,1284);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1285_up.packet_count,1285);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1286_up.packet_count,1286);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1287_up.packet_count,1287);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1288_up.packet_count,1288);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1289_up.packet_count,1289);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1290_up.packet_count,1290);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1291_up.packet_count,1291);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1292_up.packet_count,1292);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1293_up.packet_count,1293);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1294_up.packet_count,1294);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1295_up.packet_count,1295);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1296_up.packet_count,1296);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1297_up.packet_count,1297);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1298_up.packet_count,1298);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1299_up.packet_count,1299);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1300_up.packet_count,1300);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1301_up.packet_count,1301);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1302_up.packet_count,1302);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1303_up.packet_count,1303);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1304_up.packet_count,1304);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1305_up.packet_count,1305);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1306_up.packet_count,1306);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1307_up.packet_count,1307);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1308_up.packet_count,1308);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1309_up.packet_count,1309);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1310_up.packet_count,1310);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1311_up.packet_count,1311);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1312_up.packet_count,1312);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1313_up.packet_count,1313);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1314_up.packet_count,1314);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1315_up.packet_count,1315);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1316_up.packet_count,1316);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1317_up.packet_count,1317);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1318_up.packet_count,1318);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1319_up.packet_count,1319);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1320_up.packet_count,1320);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1321_up.packet_count,1321);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1322_up.packet_count,1322);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1323_up.packet_count,1323);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1324_up.packet_count,1324);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1325_up.packet_count,1325);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1326_up.packet_count,1326);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1327_up.packet_count,1327);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1328_up.packet_count,1328);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1329_up.packet_count,1329);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1330_up.packet_count,1330);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1331_up.packet_count,1331);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1332_up.packet_count,1332);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1333_up.packet_count,1333);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1334_up.packet_count,1334);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1335_up.packet_count,1335);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1336_up.packet_count,1336);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1337_up.packet_count,1337);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1338_up.packet_count,1338);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1339_up.packet_count,1339);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1340_up.packet_count,1340);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1341_up.packet_count,1341);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1342_up.packet_count,1342);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1343_up.packet_count,1343);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1344_up.packet_count,1344);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1345_up.packet_count,1345);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1346_up.packet_count,1346);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1347_up.packet_count,1347);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1348_up.packet_count,1348);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1349_up.packet_count,1349);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1350_up.packet_count,1350);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1351_up.packet_count,1351);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1352_up.packet_count,1352);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1353_up.packet_count,1353);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1354_up.packet_count,1354);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1355_up.packet_count,1355);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1356_up.packet_count,1356);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1357_up.packet_count,1357);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1358_up.packet_count,1358);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1359_up.packet_count,1359);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1360_up.packet_count,1360);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1361_up.packet_count,1361);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1362_up.packet_count,1362);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1363_up.packet_count,1363);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1364_up.packet_count,1364);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1365_up.packet_count,1365);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1366_up.packet_count,1366);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1367_up.packet_count,1367);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1368_up.packet_count,1368);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1369_up.packet_count,1369);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1370_up.packet_count,1370);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1371_up.packet_count,1371);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1372_up.packet_count,1372);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1373_up.packet_count,1373);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1374_up.packet_count,1374);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1375_up.packet_count,1375);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1376_up.packet_count,1376);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1377_up.packet_count,1377);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1378_up.packet_count,1378);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1379_up.packet_count,1379);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1380_up.packet_count,1380);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1381_up.packet_count,1381);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1382_up.packet_count,1382);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1383_up.packet_count,1383);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1384_up.packet_count,1384);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1385_up.packet_count,1385);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1386_up.packet_count,1386);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1387_up.packet_count,1387);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1388_up.packet_count,1388);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1389_up.packet_count,1389);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1390_up.packet_count,1390);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1391_up.packet_count,1391);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1392_up.packet_count,1392);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1393_up.packet_count,1393);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1394_up.packet_count,1394);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1395_up.packet_count,1395);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1396_up.packet_count,1396);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1397_up.packet_count,1397);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1398_up.packet_count,1398);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1399_up.packet_count,1399);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1400_up.packet_count,1400);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1401_up.packet_count,1401);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1402_up.packet_count,1402);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1403_up.packet_count,1403);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1404_up.packet_count,1404);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1405_up.packet_count,1405);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1406_up.packet_count,1406);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1407_up.packet_count,1407);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1408_up.packet_count,1408);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1409_up.packet_count,1409);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1410_up.packet_count,1410);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1411_up.packet_count,1411);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1412_up.packet_count,1412);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1413_up.packet_count,1413);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1414_up.packet_count,1414);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1415_up.packet_count,1415);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1416_up.packet_count,1416);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1417_up.packet_count,1417);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1418_up.packet_count,1418);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1419_up.packet_count,1419);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1420_up.packet_count,1420);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1421_up.packet_count,1421);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1422_up.packet_count,1422);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1423_up.packet_count,1423);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1424_up.packet_count,1424);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1425_up.packet_count,1425);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1426_up.packet_count,1426);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1427_up.packet_count,1427);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1428_up.packet_count,1428);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1429_up.packet_count,1429);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1430_up.packet_count,1430);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1431_up.packet_count,1431);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1432_up.packet_count,1432);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1433_up.packet_count,1433);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1434_up.packet_count,1434);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1435_up.packet_count,1435);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1436_up.packet_count,1436);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1437_up.packet_count,1437);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1438_up.packet_count,1438);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1439_up.packet_count,1439);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1440_up.packet_count,1440);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1441_up.packet_count,1441);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1442_up.packet_count,1442);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1443_up.packet_count,1443);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1444_up.packet_count,1444);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1445_up.packet_count,1445);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1446_up.packet_count,1446);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1447_up.packet_count,1447);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1448_up.packet_count,1448);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1449_up.packet_count,1449);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1450_up.packet_count,1450);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1451_up.packet_count,1451);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1452_up.packet_count,1452);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1453_up.packet_count,1453);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1454_up.packet_count,1454);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1455_up.packet_count,1455);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1456_up.packet_count,1456);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1457_up.packet_count,1457);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1458_up.packet_count,1458);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1459_up.packet_count,1459);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1460_up.packet_count,1460);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1461_up.packet_count,1461);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1462_up.packet_count,1462);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1463_up.packet_count,1463);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1464_up.packet_count,1464);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1465_up.packet_count,1465);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1466_up.packet_count,1466);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1467_up.packet_count,1467);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1468_up.packet_count,1468);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1469_up.packet_count,1469);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1470_up.packet_count,1470);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1471_up.packet_count,1471);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1472_up.packet_count,1472);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1473_up.packet_count,1473);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1474_up.packet_count,1474);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1475_up.packet_count,1475);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1476_up.packet_count,1476);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1477_up.packet_count,1477);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1478_up.packet_count,1478);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1479_up.packet_count,1479);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1480_up.packet_count,1480);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1481_up.packet_count,1481);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1482_up.packet_count,1482);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1483_up.packet_count,1483);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1484_up.packet_count,1484);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1485_up.packet_count,1485);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1486_up.packet_count,1486);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1487_up.packet_count,1487);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1488_up.packet_count,1488);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1489_up.packet_count,1489);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1490_up.packet_count,1490);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1491_up.packet_count,1491);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1492_up.packet_count,1492);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1493_up.packet_count,1493);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1494_up.packet_count,1494);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1495_up.packet_count,1495);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1496_up.packet_count,1496);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1497_up.packet_count,1497);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1498_up.packet_count,1498);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1499_up.packet_count,1499);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1500_up.packet_count,1500);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1501_up.packet_count,1501);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1502_up.packet_count,1502);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1503_up.packet_count,1503);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1504_up.packet_count,1504);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1505_up.packet_count,1505);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1506_up.packet_count,1506);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1507_up.packet_count,1507);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1508_up.packet_count,1508);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1509_up.packet_count,1509);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1510_up.packet_count,1510);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1511_up.packet_count,1511);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1512_up.packet_count,1512);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1513_up.packet_count,1513);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1514_up.packet_count,1514);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1515_up.packet_count,1515);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1516_up.packet_count,1516);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1517_up.packet_count,1517);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1518_up.packet_count,1518);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1519_up.packet_count,1519);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1520_up.packet_count,1520);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1521_up.packet_count,1521);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1522_up.packet_count,1522);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1523_up.packet_count,1523);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1524_up.packet_count,1524);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1525_up.packet_count,1525);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1526_up.packet_count,1526);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1527_up.packet_count,1527);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1528_up.packet_count,1528);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1529_up.packet_count,1529);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1530_up.packet_count,1530);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1531_up.packet_count,1531);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1532_up.packet_count,1532);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1533_up.packet_count,1533);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1534_up.packet_count,1534);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1535_up.packet_count,1535);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1536_up.packet_count,1536);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1537_up.packet_count,1537);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1538_up.packet_count,1538);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1539_up.packet_count,1539);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1540_up.packet_count,1540);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1541_up.packet_count,1541);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1542_up.packet_count,1542);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1543_up.packet_count,1543);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1544_up.packet_count,1544);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1545_up.packet_count,1545);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1546_up.packet_count,1546);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1547_up.packet_count,1547);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1548_up.packet_count,1548);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1549_up.packet_count,1549);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1550_up.packet_count,1550);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1551_up.packet_count,1551);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1552_up.packet_count,1552);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1553_up.packet_count,1553);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1554_up.packet_count,1554);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1555_up.packet_count,1555);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1556_up.packet_count,1556);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1557_up.packet_count,1557);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1558_up.packet_count,1558);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1559_up.packet_count,1559);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1560_up.packet_count,1560);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1561_up.packet_count,1561);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1562_up.packet_count,1562);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1563_up.packet_count,1563);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1564_up.packet_count,1564);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1565_up.packet_count,1565);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1566_up.packet_count,1566);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1567_up.packet_count,1567);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1568_up.packet_count,1568);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1569_up.packet_count,1569);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1570_up.packet_count,1570);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1571_up.packet_count,1571);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1572_up.packet_count,1572);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1573_up.packet_count,1573);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1574_up.packet_count,1574);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1575_up.packet_count,1575);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1576_up.packet_count,1576);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1577_up.packet_count,1577);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1578_up.packet_count,1578);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1579_up.packet_count,1579);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1580_up.packet_count,1580);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1581_up.packet_count,1581);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1582_up.packet_count,1582);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1583_up.packet_count,1583);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1584_up.packet_count,1584);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1585_up.packet_count,1585);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1586_up.packet_count,1586);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1587_up.packet_count,1587);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1588_up.packet_count,1588);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1589_up.packet_count,1589);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1590_up.packet_count,1590);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1591_up.packet_count,1591);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1592_up.packet_count,1592);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1593_up.packet_count,1593);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1594_up.packet_count,1594);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1595_up.packet_count,1595);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1596_up.packet_count,1596);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1597_up.packet_count,1597);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1598_up.packet_count,1598);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1599_up.packet_count,1599);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1600_up.packet_count,1600);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1601_up.packet_count,1601);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1602_up.packet_count,1602);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1603_up.packet_count,1603);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1604_up.packet_count,1604);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1605_up.packet_count,1605);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1606_up.packet_count,1606);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1607_up.packet_count,1607);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1608_up.packet_count,1608);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1609_up.packet_count,1609);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1610_up.packet_count,1610);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1611_up.packet_count,1611);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1612_up.packet_count,1612);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1613_up.packet_count,1613);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1614_up.packet_count,1614);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1615_up.packet_count,1615);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1616_up.packet_count,1616);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1617_up.packet_count,1617);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1618_up.packet_count,1618);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1619_up.packet_count,1619);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1620_up.packet_count,1620);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1621_up.packet_count,1621);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1622_up.packet_count,1622);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1623_up.packet_count,1623);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1624_up.packet_count,1624);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1625_up.packet_count,1625);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1626_up.packet_count,1626);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1627_up.packet_count,1627);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1628_up.packet_count,1628);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1629_up.packet_count,1629);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1630_up.packet_count,1630);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1631_up.packet_count,1631);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1632_up.packet_count,1632);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1633_up.packet_count,1633);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1634_up.packet_count,1634);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1635_up.packet_count,1635);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1636_up.packet_count,1636);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1637_up.packet_count,1637);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1638_up.packet_count,1638);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1639_up.packet_count,1639);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1640_up.packet_count,1640);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1641_up.packet_count,1641);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1642_up.packet_count,1642);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1643_up.packet_count,1643);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1644_up.packet_count,1644);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1645_up.packet_count,1645);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1646_up.packet_count,1646);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1647_up.packet_count,1647);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1648_up.packet_count,1648);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1649_up.packet_count,1649);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1650_up.packet_count,1650);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1651_up.packet_count,1651);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1652_up.packet_count,1652);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1653_up.packet_count,1653);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1654_up.packet_count,1654);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1655_up.packet_count,1655);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1656_up.packet_count,1656);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1657_up.packet_count,1657);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1658_up.packet_count,1658);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1659_up.packet_count,1659);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1660_up.packet_count,1660);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1661_up.packet_count,1661);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1662_up.packet_count,1662);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1663_up.packet_count,1663);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1664_up.packet_count,1664);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1665_up.packet_count,1665);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1666_up.packet_count,1666);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1667_up.packet_count,1667);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1668_up.packet_count,1668);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1669_up.packet_count,1669);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1670_up.packet_count,1670);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1671_up.packet_count,1671);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1672_up.packet_count,1672);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1673_up.packet_count,1673);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1674_up.packet_count,1674);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1675_up.packet_count,1675);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1676_up.packet_count,1676);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1677_up.packet_count,1677);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1678_up.packet_count,1678);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1679_up.packet_count,1679);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1680_up.packet_count,1680);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1681_up.packet_count,1681);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1682_up.packet_count,1682);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1683_up.packet_count,1683);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1684_up.packet_count,1684);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1685_up.packet_count,1685);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1686_up.packet_count,1686);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1687_up.packet_count,1687);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1688_up.packet_count,1688);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1689_up.packet_count,1689);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1690_up.packet_count,1690);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1691_up.packet_count,1691);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1692_up.packet_count,1692);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1693_up.packet_count,1693);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1694_up.packet_count,1694);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1695_up.packet_count,1695);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1696_up.packet_count,1696);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1697_up.packet_count,1697);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1698_up.packet_count,1698);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1699_up.packet_count,1699);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1700_up.packet_count,1700);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1701_up.packet_count,1701);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1702_up.packet_count,1702);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1703_up.packet_count,1703);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1704_up.packet_count,1704);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1705_up.packet_count,1705);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1706_up.packet_count,1706);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1707_up.packet_count,1707);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1708_up.packet_count,1708);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1709_up.packet_count,1709);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1710_up.packet_count,1710);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1711_up.packet_count,1711);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1712_up.packet_count,1712);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1713_up.packet_count,1713);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1714_up.packet_count,1714);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1715_up.packet_count,1715);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1716_up.packet_count,1716);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1717_up.packet_count,1717);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1718_up.packet_count,1718);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1719_up.packet_count,1719);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1720_up.packet_count,1720);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1721_up.packet_count,1721);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1722_up.packet_count,1722);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1723_up.packet_count,1723);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1724_up.packet_count,1724);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1725_up.packet_count,1725);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1726_up.packet_count,1726);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1727_up.packet_count,1727);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1728_up.packet_count,1728);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1729_up.packet_count,1729);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1730_up.packet_count,1730);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1731_up.packet_count,1731);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1732_up.packet_count,1732);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1733_up.packet_count,1733);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1734_up.packet_count,1734);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1735_up.packet_count,1735);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1736_up.packet_count,1736);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1737_up.packet_count,1737);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1738_up.packet_count,1738);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1739_up.packet_count,1739);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1740_up.packet_count,1740);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1741_up.packet_count,1741);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1742_up.packet_count,1742);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1743_up.packet_count,1743);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1744_up.packet_count,1744);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1745_up.packet_count,1745);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1746_up.packet_count,1746);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1747_up.packet_count,1747);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1748_up.packet_count,1748);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1749_up.packet_count,1749);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1750_up.packet_count,1750);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1751_up.packet_count,1751);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1752_up.packet_count,1752);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1753_up.packet_count,1753);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1754_up.packet_count,1754);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1755_up.packet_count,1755);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1756_up.packet_count,1756);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1757_up.packet_count,1757);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1758_up.packet_count,1758);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1759_up.packet_count,1759);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1760_up.packet_count,1760);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1761_up.packet_count,1761);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1762_up.packet_count,1762);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1763_up.packet_count,1763);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1764_up.packet_count,1764);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1765_up.packet_count,1765);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1766_up.packet_count,1766);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1767_up.packet_count,1767);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1768_up.packet_count,1768);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1769_up.packet_count,1769);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1770_up.packet_count,1770);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1771_up.packet_count,1771);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1772_up.packet_count,1772);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1773_up.packet_count,1773);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1774_up.packet_count,1774);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1775_up.packet_count,1775);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1776_up.packet_count,1776);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1777_up.packet_count,1777);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1778_up.packet_count,1778);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1779_up.packet_count,1779);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1780_up.packet_count,1780);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1781_up.packet_count,1781);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1782_up.packet_count,1782);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1783_up.packet_count,1783);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1784_up.packet_count,1784);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1785_up.packet_count,1785);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1786_up.packet_count,1786);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1787_up.packet_count,1787);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1788_up.packet_count,1788);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1789_up.packet_count,1789);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1790_up.packet_count,1790);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1791_up.packet_count,1791);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1792_up.packet_count,1792);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1793_up.packet_count,1793);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1794_up.packet_count,1794);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1795_up.packet_count,1795);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1796_up.packet_count,1796);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1797_up.packet_count,1797);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1798_up.packet_count,1798);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1799_up.packet_count,1799);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1800_up.packet_count,1800);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1801_up.packet_count,1801);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1802_up.packet_count,1802);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1803_up.packet_count,1803);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1804_up.packet_count,1804);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1805_up.packet_count,1805);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1806_up.packet_count,1806);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1807_up.packet_count,1807);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1808_up.packet_count,1808);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1809_up.packet_count,1809);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1810_up.packet_count,1810);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1811_up.packet_count,1811);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1812_up.packet_count,1812);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1813_up.packet_count,1813);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1814_up.packet_count,1814);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1815_up.packet_count,1815);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1816_up.packet_count,1816);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1817_up.packet_count,1817);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1818_up.packet_count,1818);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1819_up.packet_count,1819);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1820_up.packet_count,1820);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1821_up.packet_count,1821);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1822_up.packet_count,1822);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1823_up.packet_count,1823);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1824_up.packet_count,1824);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1825_up.packet_count,1825);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1826_up.packet_count,1826);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1827_up.packet_count,1827);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1828_up.packet_count,1828);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1829_up.packet_count,1829);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1830_up.packet_count,1830);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1831_up.packet_count,1831);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1832_up.packet_count,1832);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1833_up.packet_count,1833);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1834_up.packet_count,1834);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1835_up.packet_count,1835);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1836_up.packet_count,1836);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1837_up.packet_count,1837);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1838_up.packet_count,1838);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1839_up.packet_count,1839);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1840_up.packet_count,1840);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1841_up.packet_count,1841);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1842_up.packet_count,1842);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1843_up.packet_count,1843);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1844_up.packet_count,1844);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1845_up.packet_count,1845);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1846_up.packet_count,1846);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1847_up.packet_count,1847);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1848_up.packet_count,1848);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1849_up.packet_count,1849);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1850_up.packet_count,1850);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1851_up.packet_count,1851);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1852_up.packet_count,1852);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1853_up.packet_count,1853);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1854_up.packet_count,1854);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1855_up.packet_count,1855);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1856_up.packet_count,1856);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1857_up.packet_count,1857);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1858_up.packet_count,1858);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1859_up.packet_count,1859);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1860_up.packet_count,1860);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1861_up.packet_count,1861);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1862_up.packet_count,1862);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1863_up.packet_count,1863);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1864_up.packet_count,1864);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1865_up.packet_count,1865);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1866_up.packet_count,1866);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1867_up.packet_count,1867);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1868_up.packet_count,1868);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1869_up.packet_count,1869);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1870_up.packet_count,1870);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1871_up.packet_count,1871);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1872_up.packet_count,1872);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1873_up.packet_count,1873);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1874_up.packet_count,1874);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1875_up.packet_count,1875);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1876_up.packet_count,1876);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1877_up.packet_count,1877);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1878_up.packet_count,1878);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1879_up.packet_count,1879);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1880_up.packet_count,1880);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1881_up.packet_count,1881);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1882_up.packet_count,1882);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1883_up.packet_count,1883);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1884_up.packet_count,1884);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1885_up.packet_count,1885);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1886_up.packet_count,1886);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1887_up.packet_count,1887);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1888_up.packet_count,1888);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1889_up.packet_count,1889);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1890_up.packet_count,1890);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1891_up.packet_count,1891);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1892_up.packet_count,1892);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1893_up.packet_count,1893);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1894_up.packet_count,1894);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1895_up.packet_count,1895);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1896_up.packet_count,1896);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1897_up.packet_count,1897);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1898_up.packet_count,1898);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1899_up.packet_count,1899);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1900_up.packet_count,1900);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1901_up.packet_count,1901);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1902_up.packet_count,1902);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1903_up.packet_count,1903);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1904_up.packet_count,1904);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1905_up.packet_count,1905);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1906_up.packet_count,1906);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1907_up.packet_count,1907);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1908_up.packet_count,1908);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1909_up.packet_count,1909);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1910_up.packet_count,1910);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1911_up.packet_count,1911);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1912_up.packet_count,1912);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1913_up.packet_count,1913);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1914_up.packet_count,1914);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1915_up.packet_count,1915);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1916_up.packet_count,1916);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1917_up.packet_count,1917);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1918_up.packet_count,1918);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1919_up.packet_count,1919);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1920_up.packet_count,1920);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1921_up.packet_count,1921);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1922_up.packet_count,1922);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1923_up.packet_count,1923);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1924_up.packet_count,1924);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1925_up.packet_count,1925);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1926_up.packet_count,1926);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1927_up.packet_count,1927);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1928_up.packet_count,1928);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1929_up.packet_count,1929);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1930_up.packet_count,1930);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1931_up.packet_count,1931);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1932_up.packet_count,1932);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1933_up.packet_count,1933);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1934_up.packet_count,1934);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1935_up.packet_count,1935);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1936_up.packet_count,1936);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1937_up.packet_count,1937);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1938_up.packet_count,1938);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1939_up.packet_count,1939);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1940_up.packet_count,1940);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1941_up.packet_count,1941);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1942_up.packet_count,1942);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1943_up.packet_count,1943);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1944_up.packet_count,1944);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1945_up.packet_count,1945);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1946_up.packet_count,1946);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1947_up.packet_count,1947);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1948_up.packet_count,1948);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1949_up.packet_count,1949);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1950_up.packet_count,1950);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1951_up.packet_count,1951);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1952_up.packet_count,1952);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1953_up.packet_count,1953);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1954_up.packet_count,1954);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1955_up.packet_count,1955);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1956_up.packet_count,1956);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1957_up.packet_count,1957);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1958_up.packet_count,1958);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1959_up.packet_count,1959);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1960_up.packet_count,1960);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1961_up.packet_count,1961);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1962_up.packet_count,1962);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1963_up.packet_count,1963);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1964_up.packet_count,1964);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1965_up.packet_count,1965);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1966_up.packet_count,1966);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1967_up.packet_count,1967);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1968_up.packet_count,1968);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1969_up.packet_count,1969);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1970_up.packet_count,1970);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1971_up.packet_count,1971);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1972_up.packet_count,1972);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1973_up.packet_count,1973);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1974_up.packet_count,1974);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1975_up.packet_count,1975);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1976_up.packet_count,1976);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1977_up.packet_count,1977);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1978_up.packet_count,1978);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1979_up.packet_count,1979);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1980_up.packet_count,1980);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1981_up.packet_count,1981);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1982_up.packet_count,1982);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1983_up.packet_count,1983);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1984_up.packet_count,1984);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1985_up.packet_count,1985);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1986_up.packet_count,1986);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1987_up.packet_count,1987);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1988_up.packet_count,1988);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1989_up.packet_count,1989);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1990_up.packet_count,1990);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1991_up.packet_count,1991);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1992_up.packet_count,1992);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1993_up.packet_count,1993);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1994_up.packet_count,1994);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1995_up.packet_count,1995);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1996_up.packet_count,1996);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1997_up.packet_count,1997);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1998_up.packet_count,1998);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_1999_up.packet_count,1999);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2000_up.packet_count,2000);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2001_up.packet_count,2001);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2002_up.packet_count,2002);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2003_up.packet_count,2003);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2004_up.packet_count,2004);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2005_up.packet_count,2005);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2006_up.packet_count,2006);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2007_up.packet_count,2007);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2008_up.packet_count,2008);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2009_up.packet_count,2009);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2010_up.packet_count,2010);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2011_up.packet_count,2011);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2012_up.packet_count,2012);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2013_up.packet_count,2013);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2014_up.packet_count,2014);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2015_up.packet_count,2015);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2016_up.packet_count,2016);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2017_up.packet_count,2017);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2018_up.packet_count,2018);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2019_up.packet_count,2019);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2020_up.packet_count,2020);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2021_up.packet_count,2021);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2022_up.packet_count,2022);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2023_up.packet_count,2023);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2024_up.packet_count,2024);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2025_up.packet_count,2025);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2026_up.packet_count,2026);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2027_up.packet_count,2027);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2028_up.packet_count,2028);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2029_up.packet_count,2029);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2030_up.packet_count,2030);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2031_up.packet_count,2031);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2032_up.packet_count,2032);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2033_up.packet_count,2033);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2034_up.packet_count,2034);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2035_up.packet_count,2035);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2036_up.packet_count,2036);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2037_up.packet_count,2037);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2038_up.packet_count,2038);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2039_up.packet_count,2039);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2040_up.packet_count,2040);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2041_up.packet_count,2041);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2042_up.packet_count,2042);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2043_up.packet_count,2043);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2044_up.packet_count,2044);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2045_up.packet_count,2045);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2046_up.packet_count,2046);
      packet_count_check(packet_count,env.pf_vf_mux_scbd_2047_up.packet_count,2047);
      `endif
  endfunction


  function packet_count_check(int packet_sent,int packet_received,int port);
      if(packet_sent != packet_received)
				begin
             `uvm_error(get_type_name(), $sformatf("Number of packets sent at port%0d = %0d | Number of packets received at port%0d = %0d",port,packet_sent,port,packet_received));
				end
			else
				 begin
             `uvm_info(get_type_name(), $sformatf("Number of packets sent at port%0d = %0d | Number of packets received at port%0d = %0d",port,packet_sent,port,packet_received),UVM_LOW);
				 end
  endfunction

  function port_sample_count_check();
		     uvm_config_db #(int)::get(null,"","PORT_0_COUNT",port_count[0]);
		     uvm_config_db #(int)::get(null,"","PORT_1_COUNT",port_count[1]);
		     uvm_config_db #(int)::get(null,"","PORT_2_COUNT",port_count[2]);
		     uvm_config_db #(int)::get(null,"","PORT_3_COUNT",port_count[3]);
		     uvm_config_db #(int)::get(null,"","PORT_4_COUNT",port_count[4]);
		     uvm_config_db #(int)::get(null,"","PORT_5_COUNT",port_count[5]);
		     uvm_config_db #(int)::get(null,"","PORT_6_COUNT",port_count[6]);
		     uvm_config_db #(int)::get(null,"","PORT_7_COUNT",port_count[7]);
		     uvm_config_db #(int)::get(null,"","PORT_8_COUNT",port_count[8]);
		     uvm_config_db #(int)::get(null,"","PORT_9_COUNT",port_count[9]);
		     uvm_config_db #(int)::get(null,"","PORT_10_COUNT",port_count[10]);
		     uvm_config_db #(int)::get(null,"","PORT_11_COUNT",port_count[11]);
		     uvm_config_db #(int)::get(null,"","PORT_12_COUNT",port_count[12]);
		     uvm_config_db #(int)::get(null,"","PORT_13_COUNT",port_count[13]);
		     uvm_config_db #(int)::get(null,"","PORT_14_COUNT",port_count[14]);
		     uvm_config_db #(int)::get(null,"","PORT_15_COUNT",port_count[15]);
		     `ifdef TB_CONFIG_2
         uvm_config_db #(int)::get(null,"","PORT_16_COUNT",port_count[16]);
		     uvm_config_db #(int)::get(null,"","PORT_17_COUNT",port_count[17]);
		     uvm_config_db #(int)::get(null,"","PORT_18_COUNT",port_count[18]);
		     uvm_config_db #(int)::get(null,"","PORT_19_COUNT",port_count[19]);
		     uvm_config_db #(int)::get(null,"","PORT_20_COUNT",port_count[20]);
		     uvm_config_db #(int)::get(null,"","PORT_21_COUNT",port_count[21]);
		     uvm_config_db #(int)::get(null,"","PORT_22_COUNT",port_count[22]);
		     uvm_config_db #(int)::get(null,"","PORT_23_COUNT",port_count[23]);         
		     `elsif TB_CONFIG_3
         uvm_config_db #(int)::get(null,"","PORT_16_COUNT",port_count[16]);
		     uvm_config_db #(int)::get(null,"","PORT_17_COUNT",port_count[17]);
		     uvm_config_db #(int)::get(null,"","PORT_18_COUNT",port_count[18]);
		     uvm_config_db #(int)::get(null,"","PORT_19_COUNT",port_count[19]);
		     uvm_config_db #(int)::get(null,"","PORT_20_COUNT",port_count[20]);
		     uvm_config_db #(int)::get(null,"","PORT_21_COUNT",port_count[21]);
		     uvm_config_db #(int)::get(null,"","PORT_22_COUNT",port_count[22]);
		     uvm_config_db #(int)::get(null,"","PORT_23_COUNT",port_count[23]);         
         uvm_config_db #(int)::get(null,"","PORT_24_COUNT",port_count[24]);
		     uvm_config_db #(int)::get(null,"","PORT_25_COUNT",port_count[25]);
		     uvm_config_db #(int)::get(null,"","PORT_26_COUNT",port_count[26]);
		     uvm_config_db #(int)::get(null,"","PORT_27_COUNT",port_count[27]);
		     uvm_config_db #(int)::get(null,"","PORT_28_COUNT",port_count[28]);
		     uvm_config_db #(int)::get(null,"","PORT_29_COUNT",port_count[29]);
		     uvm_config_db #(int)::get(null,"","PORT_30_COUNT",port_count[30]);
		     uvm_config_db #(int)::get(null,"","PORT_31_COUNT",port_count[31]);
		     `elsif TB_CONFIG_4
		     uvm_config_db #(int)::get(null,"","PORT_16_COUNT",port_count[16]);
		     uvm_config_db #(int)::get(null,"","PORT_17_COUNT",port_count[17]);
		     uvm_config_db #(int)::get(null,"","PORT_18_COUNT",port_count[18]);
		     uvm_config_db #(int)::get(null,"","PORT_19_COUNT",port_count[19]);
		     uvm_config_db #(int)::get(null,"","PORT_20_COUNT",port_count[20]);
		     uvm_config_db #(int)::get(null,"","PORT_21_COUNT",port_count[21]);
		     uvm_config_db #(int)::get(null,"","PORT_22_COUNT",port_count[22]);
		     uvm_config_db #(int)::get(null,"","PORT_23_COUNT",port_count[23]);
		     uvm_config_db #(int)::get(null,"","PORT_24_COUNT",port_count[24]);
		     uvm_config_db #(int)::get(null,"","PORT_25_COUNT",port_count[25]);
		     uvm_config_db #(int)::get(null,"","PORT_26_COUNT",port_count[26]);
		     uvm_config_db #(int)::get(null,"","PORT_27_COUNT",port_count[27]);
		     uvm_config_db #(int)::get(null,"","PORT_28_COUNT",port_count[28]);
		     uvm_config_db #(int)::get(null,"","PORT_29_COUNT",port_count[29]);
		     uvm_config_db #(int)::get(null,"","PORT_30_COUNT",port_count[30]);
		     uvm_config_db #(int)::get(null,"","PORT_31_COUNT",port_count[31]);
		     uvm_config_db #(int)::get(null,"","PORT_32_COUNT",port_count[32]);
		     uvm_config_db #(int)::get(null,"","PORT_33_COUNT",port_count[33]);
		     uvm_config_db #(int)::get(null,"","PORT_34_COUNT",port_count[34]);
		     uvm_config_db #(int)::get(null,"","PORT_35_COUNT",port_count[35]);
		     uvm_config_db #(int)::get(null,"","PORT_36_COUNT",port_count[36]);
		     uvm_config_db #(int)::get(null,"","PORT_37_COUNT",port_count[37]);
		     uvm_config_db #(int)::get(null,"","PORT_38_COUNT",port_count[38]);
		     uvm_config_db #(int)::get(null,"","PORT_39_COUNT",port_count[39]);
		     uvm_config_db #(int)::get(null,"","PORT_40_COUNT",port_count[40]);
		     uvm_config_db #(int)::get(null,"","PORT_41_COUNT",port_count[41]);
		     uvm_config_db #(int)::get(null,"","PORT_42_COUNT",port_count[42]);
		     uvm_config_db #(int)::get(null,"","PORT_43_COUNT",port_count[43]);
		     uvm_config_db #(int)::get(null,"","PORT_44_COUNT",port_count[44]);
		     uvm_config_db #(int)::get(null,"","PORT_45_COUNT",port_count[45]);
		     uvm_config_db #(int)::get(null,"","PORT_46_COUNT",port_count[46]);
		     uvm_config_db #(int)::get(null,"","PORT_47_COUNT",port_count[47]);
		     uvm_config_db #(int)::get(null,"","PORT_48_COUNT",port_count[48]);
		     uvm_config_db #(int)::get(null,"","PORT_49_COUNT",port_count[49]);
		     uvm_config_db #(int)::get(null,"","PORT_50_COUNT",port_count[50]);
		     uvm_config_db #(int)::get(null,"","PORT_51_COUNT",port_count[51]);
		     uvm_config_db #(int)::get(null,"","PORT_52_COUNT",port_count[52]);
		     uvm_config_db #(int)::get(null,"","PORT_53_COUNT",port_count[53]);
		     uvm_config_db #(int)::get(null,"","PORT_54_COUNT",port_count[54]);
		     uvm_config_db #(int)::get(null,"","PORT_55_COUNT",port_count[55]);
		     uvm_config_db #(int)::get(null,"","PORT_56_COUNT",port_count[56]);
		     uvm_config_db #(int)::get(null,"","PORT_57_COUNT",port_count[57]);
		     uvm_config_db #(int)::get(null,"","PORT_58_COUNT",port_count[58]);
		     uvm_config_db #(int)::get(null,"","PORT_59_COUNT",port_count[59]);
		     uvm_config_db #(int)::get(null,"","PORT_60_COUNT",port_count[60]);
		     uvm_config_db #(int)::get(null,"","PORT_61_COUNT",port_count[61]);
		     uvm_config_db #(int)::get(null,"","PORT_62_COUNT",port_count[62]);
		     uvm_config_db #(int)::get(null,"","PORT_63_COUNT",port_count[63]);
		     uvm_config_db #(int)::get(null,"","PORT_64_COUNT",port_count[64]);
		     uvm_config_db #(int)::get(null,"","PORT_65_COUNT",port_count[65]);
		     uvm_config_db #(int)::get(null,"","PORT_66_COUNT",port_count[66]);
		     uvm_config_db #(int)::get(null,"","PORT_67_COUNT",port_count[67]);
		     uvm_config_db #(int)::get(null,"","PORT_68_COUNT",port_count[68]);
		     uvm_config_db #(int)::get(null,"","PORT_69_COUNT",port_count[69]);
		     uvm_config_db #(int)::get(null,"","PORT_70_COUNT",port_count[70]);
		     uvm_config_db #(int)::get(null,"","PORT_71_COUNT",port_count[71]);
		     uvm_config_db #(int)::get(null,"","PORT_72_COUNT",port_count[72]);
		     uvm_config_db #(int)::get(null,"","PORT_73_COUNT",port_count[73]);
		     uvm_config_db #(int)::get(null,"","PORT_74_COUNT",port_count[74]);
		     uvm_config_db #(int)::get(null,"","PORT_75_COUNT",port_count[75]);
		     uvm_config_db #(int)::get(null,"","PORT_76_COUNT",port_count[76]);
		     uvm_config_db #(int)::get(null,"","PORT_77_COUNT",port_count[77]);
		     uvm_config_db #(int)::get(null,"","PORT_78_COUNT",port_count[78]);
		     uvm_config_db #(int)::get(null,"","PORT_79_COUNT",port_count[79]);
		     uvm_config_db #(int)::get(null,"","PORT_80_COUNT",port_count[80]);
		     uvm_config_db #(int)::get(null,"","PORT_81_COUNT",port_count[81]);
		     uvm_config_db #(int)::get(null,"","PORT_82_COUNT",port_count[82]);
		     uvm_config_db #(int)::get(null,"","PORT_83_COUNT",port_count[83]);
		     uvm_config_db #(int)::get(null,"","PORT_84_COUNT",port_count[84]);
		     uvm_config_db #(int)::get(null,"","PORT_85_COUNT",port_count[85]);
		     uvm_config_db #(int)::get(null,"","PORT_86_COUNT",port_count[86]);
		     uvm_config_db #(int)::get(null,"","PORT_87_COUNT",port_count[87]);
		     uvm_config_db #(int)::get(null,"","PORT_88_COUNT",port_count[88]);
		     uvm_config_db #(int)::get(null,"","PORT_89_COUNT",port_count[89]);
		     uvm_config_db #(int)::get(null,"","PORT_90_COUNT",port_count[90]);
		     uvm_config_db #(int)::get(null,"","PORT_91_COUNT",port_count[91]);
		     uvm_config_db #(int)::get(null,"","PORT_92_COUNT",port_count[92]);
		     uvm_config_db #(int)::get(null,"","PORT_93_COUNT",port_count[93]);
		     uvm_config_db #(int)::get(null,"","PORT_94_COUNT",port_count[94]);
		     uvm_config_db #(int)::get(null,"","PORT_95_COUNT",port_count[95]);
		     uvm_config_db #(int)::get(null,"","PORT_96_COUNT",port_count[96]);
		     uvm_config_db #(int)::get(null,"","PORT_97_COUNT",port_count[97]);
		     uvm_config_db #(int)::get(null,"","PORT_98_COUNT",port_count[98]);
		     uvm_config_db #(int)::get(null,"","PORT_99_COUNT",port_count[99]);
		     uvm_config_db #(int)::get(null,"","PORT_100_COUNT",port_count[100]);
		     uvm_config_db #(int)::get(null,"","PORT_101_COUNT",port_count[101]);
		     uvm_config_db #(int)::get(null,"","PORT_102_COUNT",port_count[102]);
		     uvm_config_db #(int)::get(null,"","PORT_103_COUNT",port_count[103]);
		     uvm_config_db #(int)::get(null,"","PORT_104_COUNT",port_count[104]);
		     uvm_config_db #(int)::get(null,"","PORT_105_COUNT",port_count[105]);
		     uvm_config_db #(int)::get(null,"","PORT_106_COUNT",port_count[106]);
		     uvm_config_db #(int)::get(null,"","PORT_107_COUNT",port_count[107]);
		     uvm_config_db #(int)::get(null,"","PORT_108_COUNT",port_count[108]);
		     uvm_config_db #(int)::get(null,"","PORT_109_COUNT",port_count[109]);
		     uvm_config_db #(int)::get(null,"","PORT_110_COUNT",port_count[110]);
		     uvm_config_db #(int)::get(null,"","PORT_111_COUNT",port_count[111]);
		     uvm_config_db #(int)::get(null,"","PORT_112_COUNT",port_count[112]);
		     uvm_config_db #(int)::get(null,"","PORT_113_COUNT",port_count[113]);
		     uvm_config_db #(int)::get(null,"","PORT_114_COUNT",port_count[114]);
		     uvm_config_db #(int)::get(null,"","PORT_115_COUNT",port_count[115]);
		     uvm_config_db #(int)::get(null,"","PORT_116_COUNT",port_count[116]);
		     uvm_config_db #(int)::get(null,"","PORT_117_COUNT",port_count[117]);
		     uvm_config_db #(int)::get(null,"","PORT_118_COUNT",port_count[118]);
		     uvm_config_db #(int)::get(null,"","PORT_119_COUNT",port_count[119]);
		     uvm_config_db #(int)::get(null,"","PORT_120_COUNT",port_count[120]);
		     uvm_config_db #(int)::get(null,"","PORT_121_COUNT",port_count[121]);
		     uvm_config_db #(int)::get(null,"","PORT_122_COUNT",port_count[122]);
		     uvm_config_db #(int)::get(null,"","PORT_123_COUNT",port_count[123]);
		     uvm_config_db #(int)::get(null,"","PORT_124_COUNT",port_count[124]);
		     uvm_config_db #(int)::get(null,"","PORT_125_COUNT",port_count[125]);
		     uvm_config_db #(int)::get(null,"","PORT_126_COUNT",port_count[126]);
		     uvm_config_db #(int)::get(null,"","PORT_127_COUNT",port_count[127]);
		     uvm_config_db #(int)::get(null,"","PORT_128_COUNT",port_count[128]);
		     uvm_config_db #(int)::get(null,"","PORT_129_COUNT",port_count[129]);
		     uvm_config_db #(int)::get(null,"","PORT_130_COUNT",port_count[130]);
		     uvm_config_db #(int)::get(null,"","PORT_131_COUNT",port_count[131]);
		     uvm_config_db #(int)::get(null,"","PORT_132_COUNT",port_count[132]);
		     uvm_config_db #(int)::get(null,"","PORT_133_COUNT",port_count[133]);
		     uvm_config_db #(int)::get(null,"","PORT_134_COUNT",port_count[134]);
		     uvm_config_db #(int)::get(null,"","PORT_135_COUNT",port_count[135]);
		     uvm_config_db #(int)::get(null,"","PORT_136_COUNT",port_count[136]);
		     uvm_config_db #(int)::get(null,"","PORT_137_COUNT",port_count[137]);
		     uvm_config_db #(int)::get(null,"","PORT_138_COUNT",port_count[138]);
		     uvm_config_db #(int)::get(null,"","PORT_139_COUNT",port_count[139]);
		     uvm_config_db #(int)::get(null,"","PORT_140_COUNT",port_count[140]);
		     uvm_config_db #(int)::get(null,"","PORT_141_COUNT",port_count[141]);
		     uvm_config_db #(int)::get(null,"","PORT_142_COUNT",port_count[142]);
		     uvm_config_db #(int)::get(null,"","PORT_143_COUNT",port_count[143]);
		     uvm_config_db #(int)::get(null,"","PORT_144_COUNT",port_count[144]);
		     uvm_config_db #(int)::get(null,"","PORT_145_COUNT",port_count[145]);
		     uvm_config_db #(int)::get(null,"","PORT_146_COUNT",port_count[146]);
		     uvm_config_db #(int)::get(null,"","PORT_147_COUNT",port_count[147]);
		     uvm_config_db #(int)::get(null,"","PORT_148_COUNT",port_count[148]);
		     uvm_config_db #(int)::get(null,"","PORT_149_COUNT",port_count[149]);
		     uvm_config_db #(int)::get(null,"","PORT_150_COUNT",port_count[150]);
		     uvm_config_db #(int)::get(null,"","PORT_151_COUNT",port_count[151]);
		     uvm_config_db #(int)::get(null,"","PORT_152_COUNT",port_count[152]);
		     uvm_config_db #(int)::get(null,"","PORT_153_COUNT",port_count[153]);
		     uvm_config_db #(int)::get(null,"","PORT_154_COUNT",port_count[154]);
		     uvm_config_db #(int)::get(null,"","PORT_155_COUNT",port_count[155]);
		     uvm_config_db #(int)::get(null,"","PORT_156_COUNT",port_count[156]);
		     uvm_config_db #(int)::get(null,"","PORT_157_COUNT",port_count[157]);
		     uvm_config_db #(int)::get(null,"","PORT_158_COUNT",port_count[158]);
		     uvm_config_db #(int)::get(null,"","PORT_159_COUNT",port_count[159]);
		     uvm_config_db #(int)::get(null,"","PORT_160_COUNT",port_count[160]);
		     uvm_config_db #(int)::get(null,"","PORT_161_COUNT",port_count[161]);
		     uvm_config_db #(int)::get(null,"","PORT_162_COUNT",port_count[162]);
		     uvm_config_db #(int)::get(null,"","PORT_163_COUNT",port_count[163]);
		     uvm_config_db #(int)::get(null,"","PORT_164_COUNT",port_count[164]);
		     uvm_config_db #(int)::get(null,"","PORT_165_COUNT",port_count[165]);
		     uvm_config_db #(int)::get(null,"","PORT_166_COUNT",port_count[166]);
		     uvm_config_db #(int)::get(null,"","PORT_167_COUNT",port_count[167]);
		     uvm_config_db #(int)::get(null,"","PORT_168_COUNT",port_count[168]);
		     uvm_config_db #(int)::get(null,"","PORT_169_COUNT",port_count[169]);
		     uvm_config_db #(int)::get(null,"","PORT_170_COUNT",port_count[170]);
		     uvm_config_db #(int)::get(null,"","PORT_171_COUNT",port_count[171]);
		     uvm_config_db #(int)::get(null,"","PORT_172_COUNT",port_count[172]);
		     uvm_config_db #(int)::get(null,"","PORT_173_COUNT",port_count[173]);
		     uvm_config_db #(int)::get(null,"","PORT_174_COUNT",port_count[174]);
		     uvm_config_db #(int)::get(null,"","PORT_175_COUNT",port_count[175]);
		     uvm_config_db #(int)::get(null,"","PORT_176_COUNT",port_count[176]);
		     uvm_config_db #(int)::get(null,"","PORT_177_COUNT",port_count[177]);
		     uvm_config_db #(int)::get(null,"","PORT_178_COUNT",port_count[178]);
		     uvm_config_db #(int)::get(null,"","PORT_179_COUNT",port_count[179]);
		     uvm_config_db #(int)::get(null,"","PORT_180_COUNT",port_count[180]);
		     uvm_config_db #(int)::get(null,"","PORT_181_COUNT",port_count[181]);
		     uvm_config_db #(int)::get(null,"","PORT_182_COUNT",port_count[182]);
		     uvm_config_db #(int)::get(null,"","PORT_183_COUNT",port_count[183]);
		     uvm_config_db #(int)::get(null,"","PORT_184_COUNT",port_count[184]);
		     uvm_config_db #(int)::get(null,"","PORT_185_COUNT",port_count[185]);
		     uvm_config_db #(int)::get(null,"","PORT_186_COUNT",port_count[186]);
		     uvm_config_db #(int)::get(null,"","PORT_187_COUNT",port_count[187]);
		     uvm_config_db #(int)::get(null,"","PORT_188_COUNT",port_count[188]);
		     uvm_config_db #(int)::get(null,"","PORT_189_COUNT",port_count[189]);
		     uvm_config_db #(int)::get(null,"","PORT_190_COUNT",port_count[190]);
		     uvm_config_db #(int)::get(null,"","PORT_191_COUNT",port_count[191]);
		     uvm_config_db #(int)::get(null,"","PORT_192_COUNT",port_count[192]);
		     uvm_config_db #(int)::get(null,"","PORT_193_COUNT",port_count[193]);
		     uvm_config_db #(int)::get(null,"","PORT_194_COUNT",port_count[194]);
		     uvm_config_db #(int)::get(null,"","PORT_195_COUNT",port_count[195]);
		     uvm_config_db #(int)::get(null,"","PORT_196_COUNT",port_count[196]);
		     uvm_config_db #(int)::get(null,"","PORT_197_COUNT",port_count[197]);
		     uvm_config_db #(int)::get(null,"","PORT_198_COUNT",port_count[198]);
		     uvm_config_db #(int)::get(null,"","PORT_199_COUNT",port_count[199]);
		     uvm_config_db #(int)::get(null,"","PORT_200_COUNT",port_count[200]);
		     uvm_config_db #(int)::get(null,"","PORT_201_COUNT",port_count[201]);
		     uvm_config_db #(int)::get(null,"","PORT_202_COUNT",port_count[202]);
		     uvm_config_db #(int)::get(null,"","PORT_203_COUNT",port_count[203]);
		     uvm_config_db #(int)::get(null,"","PORT_204_COUNT",port_count[204]);
		     uvm_config_db #(int)::get(null,"","PORT_205_COUNT",port_count[205]);
		     uvm_config_db #(int)::get(null,"","PORT_206_COUNT",port_count[206]);
		     uvm_config_db #(int)::get(null,"","PORT_207_COUNT",port_count[207]);
		     uvm_config_db #(int)::get(null,"","PORT_208_COUNT",port_count[208]);
		     uvm_config_db #(int)::get(null,"","PORT_209_COUNT",port_count[209]);
		     uvm_config_db #(int)::get(null,"","PORT_210_COUNT",port_count[210]);
		     uvm_config_db #(int)::get(null,"","PORT_211_COUNT",port_count[211]);
		     uvm_config_db #(int)::get(null,"","PORT_212_COUNT",port_count[212]);
		     uvm_config_db #(int)::get(null,"","PORT_213_COUNT",port_count[213]);
		     uvm_config_db #(int)::get(null,"","PORT_214_COUNT",port_count[214]);
		     uvm_config_db #(int)::get(null,"","PORT_215_COUNT",port_count[215]);
		     uvm_config_db #(int)::get(null,"","PORT_216_COUNT",port_count[216]);
		     uvm_config_db #(int)::get(null,"","PORT_217_COUNT",port_count[217]);
		     uvm_config_db #(int)::get(null,"","PORT_218_COUNT",port_count[218]);
		     uvm_config_db #(int)::get(null,"","PORT_219_COUNT",port_count[219]);
		     uvm_config_db #(int)::get(null,"","PORT_220_COUNT",port_count[220]);
		     uvm_config_db #(int)::get(null,"","PORT_221_COUNT",port_count[221]);
		     uvm_config_db #(int)::get(null,"","PORT_222_COUNT",port_count[222]);
		     uvm_config_db #(int)::get(null,"","PORT_223_COUNT",port_count[223]);
		     uvm_config_db #(int)::get(null,"","PORT_224_COUNT",port_count[224]);
		     uvm_config_db #(int)::get(null,"","PORT_225_COUNT",port_count[225]);
		     uvm_config_db #(int)::get(null,"","PORT_226_COUNT",port_count[226]);
		     uvm_config_db #(int)::get(null,"","PORT_227_COUNT",port_count[227]);
		     uvm_config_db #(int)::get(null,"","PORT_228_COUNT",port_count[228]);
		     uvm_config_db #(int)::get(null,"","PORT_229_COUNT",port_count[229]);
		     uvm_config_db #(int)::get(null,"","PORT_230_COUNT",port_count[230]);
		     uvm_config_db #(int)::get(null,"","PORT_231_COUNT",port_count[231]);
		     uvm_config_db #(int)::get(null,"","PORT_232_COUNT",port_count[232]);
		     uvm_config_db #(int)::get(null,"","PORT_233_COUNT",port_count[233]);
		     uvm_config_db #(int)::get(null,"","PORT_234_COUNT",port_count[234]);
		     uvm_config_db #(int)::get(null,"","PORT_235_COUNT",port_count[235]);
		     uvm_config_db #(int)::get(null,"","PORT_236_COUNT",port_count[236]);
		     uvm_config_db #(int)::get(null,"","PORT_237_COUNT",port_count[237]);
		     uvm_config_db #(int)::get(null,"","PORT_238_COUNT",port_count[238]);
		     uvm_config_db #(int)::get(null,"","PORT_239_COUNT",port_count[239]);
		     uvm_config_db #(int)::get(null,"","PORT_240_COUNT",port_count[240]);
		     uvm_config_db #(int)::get(null,"","PORT_241_COUNT",port_count[241]);
		     uvm_config_db #(int)::get(null,"","PORT_242_COUNT",port_count[242]);
		     uvm_config_db #(int)::get(null,"","PORT_243_COUNT",port_count[243]);
		     uvm_config_db #(int)::get(null,"","PORT_244_COUNT",port_count[244]);
		     uvm_config_db #(int)::get(null,"","PORT_245_COUNT",port_count[245]);
		     uvm_config_db #(int)::get(null,"","PORT_246_COUNT",port_count[246]);
		     uvm_config_db #(int)::get(null,"","PORT_247_COUNT",port_count[247]);
		     uvm_config_db #(int)::get(null,"","PORT_248_COUNT",port_count[248]);
		     uvm_config_db #(int)::get(null,"","PORT_249_COUNT",port_count[249]);
		     uvm_config_db #(int)::get(null,"","PORT_250_COUNT",port_count[250]);
		     uvm_config_db #(int)::get(null,"","PORT_251_COUNT",port_count[251]);
		     uvm_config_db #(int)::get(null,"","PORT_252_COUNT",port_count[252]);
		     uvm_config_db #(int)::get(null,"","PORT_253_COUNT",port_count[253]);
		     uvm_config_db #(int)::get(null,"","PORT_254_COUNT",port_count[254]);
		     uvm_config_db #(int)::get(null,"","PORT_255_COUNT",port_count[255]);
		     uvm_config_db #(int)::get(null,"","PORT_256_COUNT",port_count[256]);
		     uvm_config_db #(int)::get(null,"","PORT_257_COUNT",port_count[257]);
		     uvm_config_db #(int)::get(null,"","PORT_258_COUNT",port_count[258]);
		     uvm_config_db #(int)::get(null,"","PORT_259_COUNT",port_count[259]);
		     uvm_config_db #(int)::get(null,"","PORT_260_COUNT",port_count[260]);
		     uvm_config_db #(int)::get(null,"","PORT_261_COUNT",port_count[261]);
		     uvm_config_db #(int)::get(null,"","PORT_262_COUNT",port_count[262]);
		     uvm_config_db #(int)::get(null,"","PORT_263_COUNT",port_count[263]);
		     uvm_config_db #(int)::get(null,"","PORT_264_COUNT",port_count[264]);
		     uvm_config_db #(int)::get(null,"","PORT_265_COUNT",port_count[265]);
		     uvm_config_db #(int)::get(null,"","PORT_266_COUNT",port_count[266]);
		     uvm_config_db #(int)::get(null,"","PORT_267_COUNT",port_count[267]);
		     uvm_config_db #(int)::get(null,"","PORT_268_COUNT",port_count[268]);
		     uvm_config_db #(int)::get(null,"","PORT_269_COUNT",port_count[269]);
		     uvm_config_db #(int)::get(null,"","PORT_270_COUNT",port_count[270]);
		     uvm_config_db #(int)::get(null,"","PORT_271_COUNT",port_count[271]);
		     uvm_config_db #(int)::get(null,"","PORT_272_COUNT",port_count[272]);
		     uvm_config_db #(int)::get(null,"","PORT_273_COUNT",port_count[273]);
		     uvm_config_db #(int)::get(null,"","PORT_274_COUNT",port_count[274]);
		     uvm_config_db #(int)::get(null,"","PORT_275_COUNT",port_count[275]);
		     uvm_config_db #(int)::get(null,"","PORT_276_COUNT",port_count[276]);
		     uvm_config_db #(int)::get(null,"","PORT_277_COUNT",port_count[277]);
		     uvm_config_db #(int)::get(null,"","PORT_278_COUNT",port_count[278]);
		     uvm_config_db #(int)::get(null,"","PORT_279_COUNT",port_count[279]);
		     uvm_config_db #(int)::get(null,"","PORT_280_COUNT",port_count[280]);
		     uvm_config_db #(int)::get(null,"","PORT_281_COUNT",port_count[281]);
		     uvm_config_db #(int)::get(null,"","PORT_282_COUNT",port_count[282]);
		     uvm_config_db #(int)::get(null,"","PORT_283_COUNT",port_count[283]);
		     uvm_config_db #(int)::get(null,"","PORT_284_COUNT",port_count[284]);
		     uvm_config_db #(int)::get(null,"","PORT_285_COUNT",port_count[285]);
		     uvm_config_db #(int)::get(null,"","PORT_286_COUNT",port_count[286]);
		     uvm_config_db #(int)::get(null,"","PORT_287_COUNT",port_count[287]);
		     uvm_config_db #(int)::get(null,"","PORT_288_COUNT",port_count[288]);
		     uvm_config_db #(int)::get(null,"","PORT_289_COUNT",port_count[289]);
		     uvm_config_db #(int)::get(null,"","PORT_290_COUNT",port_count[290]);
		     uvm_config_db #(int)::get(null,"","PORT_291_COUNT",port_count[291]);
		     uvm_config_db #(int)::get(null,"","PORT_292_COUNT",port_count[292]);
		     uvm_config_db #(int)::get(null,"","PORT_293_COUNT",port_count[293]);
		     uvm_config_db #(int)::get(null,"","PORT_294_COUNT",port_count[294]);
		     uvm_config_db #(int)::get(null,"","PORT_295_COUNT",port_count[295]);
		     uvm_config_db #(int)::get(null,"","PORT_296_COUNT",port_count[296]);
		     uvm_config_db #(int)::get(null,"","PORT_297_COUNT",port_count[297]);
		     uvm_config_db #(int)::get(null,"","PORT_298_COUNT",port_count[298]);
		     uvm_config_db #(int)::get(null,"","PORT_299_COUNT",port_count[299]);
		     uvm_config_db #(int)::get(null,"","PORT_300_COUNT",port_count[300]);
		     uvm_config_db #(int)::get(null,"","PORT_301_COUNT",port_count[301]);
		     uvm_config_db #(int)::get(null,"","PORT_302_COUNT",port_count[302]);
		     uvm_config_db #(int)::get(null,"","PORT_303_COUNT",port_count[303]);
		     uvm_config_db #(int)::get(null,"","PORT_304_COUNT",port_count[304]);
		     uvm_config_db #(int)::get(null,"","PORT_305_COUNT",port_count[305]);
		     uvm_config_db #(int)::get(null,"","PORT_306_COUNT",port_count[306]);
		     uvm_config_db #(int)::get(null,"","PORT_307_COUNT",port_count[307]);
		     uvm_config_db #(int)::get(null,"","PORT_308_COUNT",port_count[308]);
		     uvm_config_db #(int)::get(null,"","PORT_309_COUNT",port_count[309]);
		     uvm_config_db #(int)::get(null,"","PORT_310_COUNT",port_count[310]);
		     uvm_config_db #(int)::get(null,"","PORT_311_COUNT",port_count[311]);
		     uvm_config_db #(int)::get(null,"","PORT_312_COUNT",port_count[312]);
		     uvm_config_db #(int)::get(null,"","PORT_313_COUNT",port_count[313]);
		     uvm_config_db #(int)::get(null,"","PORT_314_COUNT",port_count[314]);
		     uvm_config_db #(int)::get(null,"","PORT_315_COUNT",port_count[315]);
		     uvm_config_db #(int)::get(null,"","PORT_316_COUNT",port_count[316]);
		     uvm_config_db #(int)::get(null,"","PORT_317_COUNT",port_count[317]);
		     uvm_config_db #(int)::get(null,"","PORT_318_COUNT",port_count[318]);
		     uvm_config_db #(int)::get(null,"","PORT_319_COUNT",port_count[319]);
		     uvm_config_db #(int)::get(null,"","PORT_320_COUNT",port_count[320]);
		     uvm_config_db #(int)::get(null,"","PORT_321_COUNT",port_count[321]);
		     uvm_config_db #(int)::get(null,"","PORT_322_COUNT",port_count[322]);
		     uvm_config_db #(int)::get(null,"","PORT_323_COUNT",port_count[323]);
		     uvm_config_db #(int)::get(null,"","PORT_324_COUNT",port_count[324]);
		     uvm_config_db #(int)::get(null,"","PORT_325_COUNT",port_count[325]);
		     uvm_config_db #(int)::get(null,"","PORT_326_COUNT",port_count[326]);
		     uvm_config_db #(int)::get(null,"","PORT_327_COUNT",port_count[327]);
		     uvm_config_db #(int)::get(null,"","PORT_328_COUNT",port_count[328]);
		     uvm_config_db #(int)::get(null,"","PORT_329_COUNT",port_count[329]);
		     uvm_config_db #(int)::get(null,"","PORT_330_COUNT",port_count[330]);
		     uvm_config_db #(int)::get(null,"","PORT_331_COUNT",port_count[331]);
		     uvm_config_db #(int)::get(null,"","PORT_332_COUNT",port_count[332]);
		     uvm_config_db #(int)::get(null,"","PORT_333_COUNT",port_count[333]);
		     uvm_config_db #(int)::get(null,"","PORT_334_COUNT",port_count[334]);
		     uvm_config_db #(int)::get(null,"","PORT_335_COUNT",port_count[335]);
		     uvm_config_db #(int)::get(null,"","PORT_336_COUNT",port_count[336]);
		     uvm_config_db #(int)::get(null,"","PORT_337_COUNT",port_count[337]);
		     uvm_config_db #(int)::get(null,"","PORT_338_COUNT",port_count[338]);
		     uvm_config_db #(int)::get(null,"","PORT_339_COUNT",port_count[339]);
		     uvm_config_db #(int)::get(null,"","PORT_340_COUNT",port_count[340]);
		     uvm_config_db #(int)::get(null,"","PORT_341_COUNT",port_count[341]);
		     uvm_config_db #(int)::get(null,"","PORT_342_COUNT",port_count[342]);
		     uvm_config_db #(int)::get(null,"","PORT_343_COUNT",port_count[343]);
		     uvm_config_db #(int)::get(null,"","PORT_344_COUNT",port_count[344]);
		     uvm_config_db #(int)::get(null,"","PORT_345_COUNT",port_count[345]);
		     uvm_config_db #(int)::get(null,"","PORT_346_COUNT",port_count[346]);
		     uvm_config_db #(int)::get(null,"","PORT_347_COUNT",port_count[347]);
		     uvm_config_db #(int)::get(null,"","PORT_348_COUNT",port_count[348]);
		     uvm_config_db #(int)::get(null,"","PORT_349_COUNT",port_count[349]);
		     uvm_config_db #(int)::get(null,"","PORT_350_COUNT",port_count[350]);
		     uvm_config_db #(int)::get(null,"","PORT_351_COUNT",port_count[351]);
		     uvm_config_db #(int)::get(null,"","PORT_352_COUNT",port_count[352]);
		     uvm_config_db #(int)::get(null,"","PORT_353_COUNT",port_count[353]);
		     uvm_config_db #(int)::get(null,"","PORT_354_COUNT",port_count[354]);
		     uvm_config_db #(int)::get(null,"","PORT_355_COUNT",port_count[355]);
		     uvm_config_db #(int)::get(null,"","PORT_356_COUNT",port_count[356]);
		     uvm_config_db #(int)::get(null,"","PORT_357_COUNT",port_count[357]);
		     uvm_config_db #(int)::get(null,"","PORT_358_COUNT",port_count[358]);
		     uvm_config_db #(int)::get(null,"","PORT_359_COUNT",port_count[359]);
		     uvm_config_db #(int)::get(null,"","PORT_360_COUNT",port_count[360]);
		     uvm_config_db #(int)::get(null,"","PORT_361_COUNT",port_count[361]);
		     uvm_config_db #(int)::get(null,"","PORT_362_COUNT",port_count[362]);
		     uvm_config_db #(int)::get(null,"","PORT_363_COUNT",port_count[363]);
		     uvm_config_db #(int)::get(null,"","PORT_364_COUNT",port_count[364]);
		     uvm_config_db #(int)::get(null,"","PORT_365_COUNT",port_count[365]);
		     uvm_config_db #(int)::get(null,"","PORT_366_COUNT",port_count[366]);
		     uvm_config_db #(int)::get(null,"","PORT_367_COUNT",port_count[367]);
		     uvm_config_db #(int)::get(null,"","PORT_368_COUNT",port_count[368]);
		     uvm_config_db #(int)::get(null,"","PORT_369_COUNT",port_count[369]);
		     uvm_config_db #(int)::get(null,"","PORT_370_COUNT",port_count[370]);
		     uvm_config_db #(int)::get(null,"","PORT_371_COUNT",port_count[371]);
		     uvm_config_db #(int)::get(null,"","PORT_372_COUNT",port_count[372]);
		     uvm_config_db #(int)::get(null,"","PORT_373_COUNT",port_count[373]);
		     uvm_config_db #(int)::get(null,"","PORT_374_COUNT",port_count[374]);
		     uvm_config_db #(int)::get(null,"","PORT_375_COUNT",port_count[375]);
		     uvm_config_db #(int)::get(null,"","PORT_376_COUNT",port_count[376]);
		     uvm_config_db #(int)::get(null,"","PORT_377_COUNT",port_count[377]);
		     uvm_config_db #(int)::get(null,"","PORT_378_COUNT",port_count[378]);
		     uvm_config_db #(int)::get(null,"","PORT_379_COUNT",port_count[379]);
		     uvm_config_db #(int)::get(null,"","PORT_380_COUNT",port_count[380]);
		     uvm_config_db #(int)::get(null,"","PORT_381_COUNT",port_count[381]);
		     uvm_config_db #(int)::get(null,"","PORT_382_COUNT",port_count[382]);
		     uvm_config_db #(int)::get(null,"","PORT_383_COUNT",port_count[383]);
		     uvm_config_db #(int)::get(null,"","PORT_384_COUNT",port_count[384]);
		     uvm_config_db #(int)::get(null,"","PORT_385_COUNT",port_count[385]);
		     uvm_config_db #(int)::get(null,"","PORT_386_COUNT",port_count[386]);
		     uvm_config_db #(int)::get(null,"","PORT_387_COUNT",port_count[387]);
		     uvm_config_db #(int)::get(null,"","PORT_388_COUNT",port_count[388]);
		     uvm_config_db #(int)::get(null,"","PORT_389_COUNT",port_count[389]);
		     uvm_config_db #(int)::get(null,"","PORT_390_COUNT",port_count[390]);
		     uvm_config_db #(int)::get(null,"","PORT_391_COUNT",port_count[391]);
		     uvm_config_db #(int)::get(null,"","PORT_392_COUNT",port_count[392]);
		     uvm_config_db #(int)::get(null,"","PORT_393_COUNT",port_count[393]);
		     uvm_config_db #(int)::get(null,"","PORT_394_COUNT",port_count[394]);
		     uvm_config_db #(int)::get(null,"","PORT_395_COUNT",port_count[395]);
		     uvm_config_db #(int)::get(null,"","PORT_396_COUNT",port_count[396]);
		     uvm_config_db #(int)::get(null,"","PORT_397_COUNT",port_count[397]);
		     uvm_config_db #(int)::get(null,"","PORT_398_COUNT",port_count[398]);
		     uvm_config_db #(int)::get(null,"","PORT_399_COUNT",port_count[399]);
		     uvm_config_db #(int)::get(null,"","PORT_400_COUNT",port_count[400]);
		     uvm_config_db #(int)::get(null,"","PORT_401_COUNT",port_count[401]);
		     uvm_config_db #(int)::get(null,"","PORT_402_COUNT",port_count[402]);
		     uvm_config_db #(int)::get(null,"","PORT_403_COUNT",port_count[403]);
		     uvm_config_db #(int)::get(null,"","PORT_404_COUNT",port_count[404]);
		     uvm_config_db #(int)::get(null,"","PORT_405_COUNT",port_count[405]);
		     uvm_config_db #(int)::get(null,"","PORT_406_COUNT",port_count[406]);
		     uvm_config_db #(int)::get(null,"","PORT_407_COUNT",port_count[407]);
		     uvm_config_db #(int)::get(null,"","PORT_408_COUNT",port_count[408]);
		     uvm_config_db #(int)::get(null,"","PORT_409_COUNT",port_count[409]);
		     uvm_config_db #(int)::get(null,"","PORT_410_COUNT",port_count[410]);
		     uvm_config_db #(int)::get(null,"","PORT_411_COUNT",port_count[411]);
		     uvm_config_db #(int)::get(null,"","PORT_412_COUNT",port_count[412]);
		     uvm_config_db #(int)::get(null,"","PORT_413_COUNT",port_count[413]);
		     uvm_config_db #(int)::get(null,"","PORT_414_COUNT",port_count[414]);
		     uvm_config_db #(int)::get(null,"","PORT_415_COUNT",port_count[415]);
		     uvm_config_db #(int)::get(null,"","PORT_416_COUNT",port_count[416]);
		     uvm_config_db #(int)::get(null,"","PORT_417_COUNT",port_count[417]);
		     uvm_config_db #(int)::get(null,"","PORT_418_COUNT",port_count[418]);
		     uvm_config_db #(int)::get(null,"","PORT_419_COUNT",port_count[419]);
		     uvm_config_db #(int)::get(null,"","PORT_420_COUNT",port_count[420]);
		     uvm_config_db #(int)::get(null,"","PORT_421_COUNT",port_count[421]);
		     uvm_config_db #(int)::get(null,"","PORT_422_COUNT",port_count[422]);
		     uvm_config_db #(int)::get(null,"","PORT_423_COUNT",port_count[423]);
		     uvm_config_db #(int)::get(null,"","PORT_424_COUNT",port_count[424]);
		     uvm_config_db #(int)::get(null,"","PORT_425_COUNT",port_count[425]);
		     uvm_config_db #(int)::get(null,"","PORT_426_COUNT",port_count[426]);
		     uvm_config_db #(int)::get(null,"","PORT_427_COUNT",port_count[427]);
		     uvm_config_db #(int)::get(null,"","PORT_428_COUNT",port_count[428]);
		     uvm_config_db #(int)::get(null,"","PORT_429_COUNT",port_count[429]);
		     uvm_config_db #(int)::get(null,"","PORT_430_COUNT",port_count[430]);
		     uvm_config_db #(int)::get(null,"","PORT_431_COUNT",port_count[431]);
		     uvm_config_db #(int)::get(null,"","PORT_432_COUNT",port_count[432]);
		     uvm_config_db #(int)::get(null,"","PORT_433_COUNT",port_count[433]);
		     uvm_config_db #(int)::get(null,"","PORT_434_COUNT",port_count[434]);
		     uvm_config_db #(int)::get(null,"","PORT_435_COUNT",port_count[435]);
		     uvm_config_db #(int)::get(null,"","PORT_436_COUNT",port_count[436]);
		     uvm_config_db #(int)::get(null,"","PORT_437_COUNT",port_count[437]);
		     uvm_config_db #(int)::get(null,"","PORT_438_COUNT",port_count[438]);
		     uvm_config_db #(int)::get(null,"","PORT_439_COUNT",port_count[439]);
		     uvm_config_db #(int)::get(null,"","PORT_440_COUNT",port_count[440]);
		     uvm_config_db #(int)::get(null,"","PORT_441_COUNT",port_count[441]);
		     uvm_config_db #(int)::get(null,"","PORT_442_COUNT",port_count[442]);
		     uvm_config_db #(int)::get(null,"","PORT_443_COUNT",port_count[443]);
		     uvm_config_db #(int)::get(null,"","PORT_444_COUNT",port_count[444]);
		     uvm_config_db #(int)::get(null,"","PORT_445_COUNT",port_count[445]);
		     uvm_config_db #(int)::get(null,"","PORT_446_COUNT",port_count[446]);
		     uvm_config_db #(int)::get(null,"","PORT_447_COUNT",port_count[447]);
		     uvm_config_db #(int)::get(null,"","PORT_448_COUNT",port_count[448]);
		     uvm_config_db #(int)::get(null,"","PORT_449_COUNT",port_count[449]);
		     uvm_config_db #(int)::get(null,"","PORT_450_COUNT",port_count[450]);
		     uvm_config_db #(int)::get(null,"","PORT_451_COUNT",port_count[451]);
		     uvm_config_db #(int)::get(null,"","PORT_452_COUNT",port_count[452]);
		     uvm_config_db #(int)::get(null,"","PORT_453_COUNT",port_count[453]);
		     uvm_config_db #(int)::get(null,"","PORT_454_COUNT",port_count[454]);
		     uvm_config_db #(int)::get(null,"","PORT_455_COUNT",port_count[455]);
		     uvm_config_db #(int)::get(null,"","PORT_456_COUNT",port_count[456]);
		     uvm_config_db #(int)::get(null,"","PORT_457_COUNT",port_count[457]);
		     uvm_config_db #(int)::get(null,"","PORT_458_COUNT",port_count[458]);
		     uvm_config_db #(int)::get(null,"","PORT_459_COUNT",port_count[459]);
		     uvm_config_db #(int)::get(null,"","PORT_460_COUNT",port_count[460]);
		     uvm_config_db #(int)::get(null,"","PORT_461_COUNT",port_count[461]);
		     uvm_config_db #(int)::get(null,"","PORT_462_COUNT",port_count[462]);
		     uvm_config_db #(int)::get(null,"","PORT_463_COUNT",port_count[463]);
		     uvm_config_db #(int)::get(null,"","PORT_464_COUNT",port_count[464]);
		     uvm_config_db #(int)::get(null,"","PORT_465_COUNT",port_count[465]);
		     uvm_config_db #(int)::get(null,"","PORT_466_COUNT",port_count[466]);
		     uvm_config_db #(int)::get(null,"","PORT_467_COUNT",port_count[467]);
		     uvm_config_db #(int)::get(null,"","PORT_468_COUNT",port_count[468]);
		     uvm_config_db #(int)::get(null,"","PORT_469_COUNT",port_count[469]);
		     uvm_config_db #(int)::get(null,"","PORT_470_COUNT",port_count[470]);
		     uvm_config_db #(int)::get(null,"","PORT_471_COUNT",port_count[471]);
		     uvm_config_db #(int)::get(null,"","PORT_472_COUNT",port_count[472]);
		     uvm_config_db #(int)::get(null,"","PORT_473_COUNT",port_count[473]);
		     uvm_config_db #(int)::get(null,"","PORT_474_COUNT",port_count[474]);
		     uvm_config_db #(int)::get(null,"","PORT_475_COUNT",port_count[475]);
		     uvm_config_db #(int)::get(null,"","PORT_476_COUNT",port_count[476]);
		     uvm_config_db #(int)::get(null,"","PORT_477_COUNT",port_count[477]);
		     uvm_config_db #(int)::get(null,"","PORT_478_COUNT",port_count[478]);
		     uvm_config_db #(int)::get(null,"","PORT_479_COUNT",port_count[479]);
		     uvm_config_db #(int)::get(null,"","PORT_480_COUNT",port_count[480]);
		     uvm_config_db #(int)::get(null,"","PORT_481_COUNT",port_count[481]);
		     uvm_config_db #(int)::get(null,"","PORT_482_COUNT",port_count[482]);
		     uvm_config_db #(int)::get(null,"","PORT_483_COUNT",port_count[483]);
		     uvm_config_db #(int)::get(null,"","PORT_484_COUNT",port_count[484]);
		     uvm_config_db #(int)::get(null,"","PORT_485_COUNT",port_count[485]);
		     uvm_config_db #(int)::get(null,"","PORT_486_COUNT",port_count[486]);
		     uvm_config_db #(int)::get(null,"","PORT_487_COUNT",port_count[487]);
		     uvm_config_db #(int)::get(null,"","PORT_488_COUNT",port_count[488]);
		     uvm_config_db #(int)::get(null,"","PORT_489_COUNT",port_count[489]);
		     uvm_config_db #(int)::get(null,"","PORT_490_COUNT",port_count[490]);
		     uvm_config_db #(int)::get(null,"","PORT_491_COUNT",port_count[491]);
		     uvm_config_db #(int)::get(null,"","PORT_492_COUNT",port_count[492]);
		     uvm_config_db #(int)::get(null,"","PORT_493_COUNT",port_count[493]);
		     uvm_config_db #(int)::get(null,"","PORT_494_COUNT",port_count[494]);
		     uvm_config_db #(int)::get(null,"","PORT_495_COUNT",port_count[495]);
		     uvm_config_db #(int)::get(null,"","PORT_496_COUNT",port_count[496]);
		     uvm_config_db #(int)::get(null,"","PORT_497_COUNT",port_count[497]);
		     uvm_config_db #(int)::get(null,"","PORT_498_COUNT",port_count[498]);
		     uvm_config_db #(int)::get(null,"","PORT_499_COUNT",port_count[499]);
		     uvm_config_db #(int)::get(null,"","PORT_500_COUNT",port_count[500]);
		     uvm_config_db #(int)::get(null,"","PORT_501_COUNT",port_count[501]);
		     uvm_config_db #(int)::get(null,"","PORT_502_COUNT",port_count[502]);
		     uvm_config_db #(int)::get(null,"","PORT_503_COUNT",port_count[503]);
		     uvm_config_db #(int)::get(null,"","PORT_504_COUNT",port_count[504]);
		     uvm_config_db #(int)::get(null,"","PORT_505_COUNT",port_count[505]);
		     uvm_config_db #(int)::get(null,"","PORT_506_COUNT",port_count[506]);
		     uvm_config_db #(int)::get(null,"","PORT_507_COUNT",port_count[507]);
		     uvm_config_db #(int)::get(null,"","PORT_508_COUNT",port_count[508]);
		     uvm_config_db #(int)::get(null,"","PORT_509_COUNT",port_count[509]);
		     uvm_config_db #(int)::get(null,"","PORT_510_COUNT",port_count[510]);
		     uvm_config_db #(int)::get(null,"","PORT_511_COUNT",port_count[511]);
		     uvm_config_db #(int)::get(null,"","PORT_512_COUNT",port_count[512]);
		     uvm_config_db #(int)::get(null,"","PORT_513_COUNT",port_count[513]);
		     uvm_config_db #(int)::get(null,"","PORT_514_COUNT",port_count[514]);
		     uvm_config_db #(int)::get(null,"","PORT_515_COUNT",port_count[515]);
		     uvm_config_db #(int)::get(null,"","PORT_516_COUNT",port_count[516]);
		     uvm_config_db #(int)::get(null,"","PORT_517_COUNT",port_count[517]);
		     uvm_config_db #(int)::get(null,"","PORT_518_COUNT",port_count[518]);
		     uvm_config_db #(int)::get(null,"","PORT_519_COUNT",port_count[519]);
		     uvm_config_db #(int)::get(null,"","PORT_520_COUNT",port_count[520]);
		     uvm_config_db #(int)::get(null,"","PORT_521_COUNT",port_count[521]);
		     uvm_config_db #(int)::get(null,"","PORT_522_COUNT",port_count[522]);
		     uvm_config_db #(int)::get(null,"","PORT_523_COUNT",port_count[523]);
		     uvm_config_db #(int)::get(null,"","PORT_524_COUNT",port_count[524]);
		     uvm_config_db #(int)::get(null,"","PORT_525_COUNT",port_count[525]);
		     uvm_config_db #(int)::get(null,"","PORT_526_COUNT",port_count[526]);
		     uvm_config_db #(int)::get(null,"","PORT_527_COUNT",port_count[527]);
		     uvm_config_db #(int)::get(null,"","PORT_528_COUNT",port_count[528]);
		     uvm_config_db #(int)::get(null,"","PORT_529_COUNT",port_count[529]);
		     uvm_config_db #(int)::get(null,"","PORT_530_COUNT",port_count[530]);
		     uvm_config_db #(int)::get(null,"","PORT_531_COUNT",port_count[531]);
		     uvm_config_db #(int)::get(null,"","PORT_532_COUNT",port_count[532]);
		     uvm_config_db #(int)::get(null,"","PORT_533_COUNT",port_count[533]);
		     uvm_config_db #(int)::get(null,"","PORT_534_COUNT",port_count[534]);
		     uvm_config_db #(int)::get(null,"","PORT_535_COUNT",port_count[535]);
		     uvm_config_db #(int)::get(null,"","PORT_536_COUNT",port_count[536]);
		     uvm_config_db #(int)::get(null,"","PORT_537_COUNT",port_count[537]);
		     uvm_config_db #(int)::get(null,"","PORT_538_COUNT",port_count[538]);
		     uvm_config_db #(int)::get(null,"","PORT_539_COUNT",port_count[539]);
		     uvm_config_db #(int)::get(null,"","PORT_540_COUNT",port_count[540]);
		     uvm_config_db #(int)::get(null,"","PORT_541_COUNT",port_count[541]);
		     uvm_config_db #(int)::get(null,"","PORT_542_COUNT",port_count[542]);
		     uvm_config_db #(int)::get(null,"","PORT_543_COUNT",port_count[543]);
		     uvm_config_db #(int)::get(null,"","PORT_544_COUNT",port_count[544]);
		     uvm_config_db #(int)::get(null,"","PORT_545_COUNT",port_count[545]);
		     uvm_config_db #(int)::get(null,"","PORT_546_COUNT",port_count[546]);
		     uvm_config_db #(int)::get(null,"","PORT_547_COUNT",port_count[547]);
		     uvm_config_db #(int)::get(null,"","PORT_548_COUNT",port_count[548]);
		     uvm_config_db #(int)::get(null,"","PORT_549_COUNT",port_count[549]);
		     uvm_config_db #(int)::get(null,"","PORT_550_COUNT",port_count[550]);
		     uvm_config_db #(int)::get(null,"","PORT_551_COUNT",port_count[551]);
		     uvm_config_db #(int)::get(null,"","PORT_552_COUNT",port_count[552]);
		     uvm_config_db #(int)::get(null,"","PORT_553_COUNT",port_count[553]);
		     uvm_config_db #(int)::get(null,"","PORT_554_COUNT",port_count[554]);
		     uvm_config_db #(int)::get(null,"","PORT_555_COUNT",port_count[555]);
		     uvm_config_db #(int)::get(null,"","PORT_556_COUNT",port_count[556]);
		     uvm_config_db #(int)::get(null,"","PORT_557_COUNT",port_count[557]);
		     uvm_config_db #(int)::get(null,"","PORT_558_COUNT",port_count[558]);
		     uvm_config_db #(int)::get(null,"","PORT_559_COUNT",port_count[559]);
		     uvm_config_db #(int)::get(null,"","PORT_560_COUNT",port_count[560]);
		     uvm_config_db #(int)::get(null,"","PORT_561_COUNT",port_count[561]);
		     uvm_config_db #(int)::get(null,"","PORT_562_COUNT",port_count[562]);
		     uvm_config_db #(int)::get(null,"","PORT_563_COUNT",port_count[563]);
		     uvm_config_db #(int)::get(null,"","PORT_564_COUNT",port_count[564]);
		     uvm_config_db #(int)::get(null,"","PORT_565_COUNT",port_count[565]);
		     uvm_config_db #(int)::get(null,"","PORT_566_COUNT",port_count[566]);
		     uvm_config_db #(int)::get(null,"","PORT_567_COUNT",port_count[567]);
		     uvm_config_db #(int)::get(null,"","PORT_568_COUNT",port_count[568]);
		     uvm_config_db #(int)::get(null,"","PORT_569_COUNT",port_count[569]);
		     uvm_config_db #(int)::get(null,"","PORT_570_COUNT",port_count[570]);
		     uvm_config_db #(int)::get(null,"","PORT_571_COUNT",port_count[571]);
		     uvm_config_db #(int)::get(null,"","PORT_572_COUNT",port_count[572]);
		     uvm_config_db #(int)::get(null,"","PORT_573_COUNT",port_count[573]);
		     uvm_config_db #(int)::get(null,"","PORT_574_COUNT",port_count[574]);
		     uvm_config_db #(int)::get(null,"","PORT_575_COUNT",port_count[575]);
		     uvm_config_db #(int)::get(null,"","PORT_576_COUNT",port_count[576]);
		     uvm_config_db #(int)::get(null,"","PORT_577_COUNT",port_count[577]);
		     uvm_config_db #(int)::get(null,"","PORT_578_COUNT",port_count[578]);
		     uvm_config_db #(int)::get(null,"","PORT_579_COUNT",port_count[579]);
		     uvm_config_db #(int)::get(null,"","PORT_580_COUNT",port_count[580]);
		     uvm_config_db #(int)::get(null,"","PORT_581_COUNT",port_count[581]);
		     uvm_config_db #(int)::get(null,"","PORT_582_COUNT",port_count[582]);
		     uvm_config_db #(int)::get(null,"","PORT_583_COUNT",port_count[583]);
		     uvm_config_db #(int)::get(null,"","PORT_584_COUNT",port_count[584]);
		     uvm_config_db #(int)::get(null,"","PORT_585_COUNT",port_count[585]);
		     uvm_config_db #(int)::get(null,"","PORT_586_COUNT",port_count[586]);
		     uvm_config_db #(int)::get(null,"","PORT_587_COUNT",port_count[587]);
		     uvm_config_db #(int)::get(null,"","PORT_588_COUNT",port_count[588]);
		     uvm_config_db #(int)::get(null,"","PORT_589_COUNT",port_count[589]);
		     uvm_config_db #(int)::get(null,"","PORT_590_COUNT",port_count[590]);
		     uvm_config_db #(int)::get(null,"","PORT_591_COUNT",port_count[591]);
		     uvm_config_db #(int)::get(null,"","PORT_592_COUNT",port_count[592]);
		     uvm_config_db #(int)::get(null,"","PORT_593_COUNT",port_count[593]);
		     uvm_config_db #(int)::get(null,"","PORT_594_COUNT",port_count[594]);
		     uvm_config_db #(int)::get(null,"","PORT_595_COUNT",port_count[595]);
		     uvm_config_db #(int)::get(null,"","PORT_596_COUNT",port_count[596]);
		     uvm_config_db #(int)::get(null,"","PORT_597_COUNT",port_count[597]);
		     uvm_config_db #(int)::get(null,"","PORT_598_COUNT",port_count[598]);
		     uvm_config_db #(int)::get(null,"","PORT_599_COUNT",port_count[599]);
		     uvm_config_db #(int)::get(null,"","PORT_600_COUNT",port_count[600]);
		     uvm_config_db #(int)::get(null,"","PORT_601_COUNT",port_count[601]);
		     uvm_config_db #(int)::get(null,"","PORT_602_COUNT",port_count[602]);
		     uvm_config_db #(int)::get(null,"","PORT_603_COUNT",port_count[603]);
		     uvm_config_db #(int)::get(null,"","PORT_604_COUNT",port_count[604]);
		     uvm_config_db #(int)::get(null,"","PORT_605_COUNT",port_count[605]);
		     uvm_config_db #(int)::get(null,"","PORT_606_COUNT",port_count[606]);
		     uvm_config_db #(int)::get(null,"","PORT_607_COUNT",port_count[607]);
		     uvm_config_db #(int)::get(null,"","PORT_608_COUNT",port_count[608]);
		     uvm_config_db #(int)::get(null,"","PORT_609_COUNT",port_count[609]);
		     uvm_config_db #(int)::get(null,"","PORT_610_COUNT",port_count[610]);
		     uvm_config_db #(int)::get(null,"","PORT_611_COUNT",port_count[611]);
		     uvm_config_db #(int)::get(null,"","PORT_612_COUNT",port_count[612]);
		     uvm_config_db #(int)::get(null,"","PORT_613_COUNT",port_count[613]);
		     uvm_config_db #(int)::get(null,"","PORT_614_COUNT",port_count[614]);
		     uvm_config_db #(int)::get(null,"","PORT_615_COUNT",port_count[615]);
		     uvm_config_db #(int)::get(null,"","PORT_616_COUNT",port_count[616]);
		     uvm_config_db #(int)::get(null,"","PORT_617_COUNT",port_count[617]);
		     uvm_config_db #(int)::get(null,"","PORT_618_COUNT",port_count[618]);
		     uvm_config_db #(int)::get(null,"","PORT_619_COUNT",port_count[619]);
		     uvm_config_db #(int)::get(null,"","PORT_620_COUNT",port_count[620]);
		     uvm_config_db #(int)::get(null,"","PORT_621_COUNT",port_count[621]);
		     uvm_config_db #(int)::get(null,"","PORT_622_COUNT",port_count[622]);
		     uvm_config_db #(int)::get(null,"","PORT_623_COUNT",port_count[623]);
		     uvm_config_db #(int)::get(null,"","PORT_624_COUNT",port_count[624]);
		     uvm_config_db #(int)::get(null,"","PORT_625_COUNT",port_count[625]);
		     uvm_config_db #(int)::get(null,"","PORT_626_COUNT",port_count[626]);
		     uvm_config_db #(int)::get(null,"","PORT_627_COUNT",port_count[627]);
		     uvm_config_db #(int)::get(null,"","PORT_628_COUNT",port_count[628]);
		     uvm_config_db #(int)::get(null,"","PORT_629_COUNT",port_count[629]);
		     uvm_config_db #(int)::get(null,"","PORT_630_COUNT",port_count[630]);
		     uvm_config_db #(int)::get(null,"","PORT_631_COUNT",port_count[631]);
		     uvm_config_db #(int)::get(null,"","PORT_632_COUNT",port_count[632]);
		     uvm_config_db #(int)::get(null,"","PORT_633_COUNT",port_count[633]);
		     uvm_config_db #(int)::get(null,"","PORT_634_COUNT",port_count[634]);
		     uvm_config_db #(int)::get(null,"","PORT_635_COUNT",port_count[635]);
		     uvm_config_db #(int)::get(null,"","PORT_636_COUNT",port_count[636]);
		     uvm_config_db #(int)::get(null,"","PORT_637_COUNT",port_count[637]);
		     uvm_config_db #(int)::get(null,"","PORT_638_COUNT",port_count[638]);
		     uvm_config_db #(int)::get(null,"","PORT_639_COUNT",port_count[639]);
		     uvm_config_db #(int)::get(null,"","PORT_640_COUNT",port_count[640]);
		     uvm_config_db #(int)::get(null,"","PORT_641_COUNT",port_count[641]);
		     uvm_config_db #(int)::get(null,"","PORT_642_COUNT",port_count[642]);
		     uvm_config_db #(int)::get(null,"","PORT_643_COUNT",port_count[643]);
		     uvm_config_db #(int)::get(null,"","PORT_644_COUNT",port_count[644]);
		     uvm_config_db #(int)::get(null,"","PORT_645_COUNT",port_count[645]);
		     uvm_config_db #(int)::get(null,"","PORT_646_COUNT",port_count[646]);
		     uvm_config_db #(int)::get(null,"","PORT_647_COUNT",port_count[647]);
		     uvm_config_db #(int)::get(null,"","PORT_648_COUNT",port_count[648]);
		     uvm_config_db #(int)::get(null,"","PORT_649_COUNT",port_count[649]);
		     uvm_config_db #(int)::get(null,"","PORT_650_COUNT",port_count[650]);
		     uvm_config_db #(int)::get(null,"","PORT_651_COUNT",port_count[651]);
		     uvm_config_db #(int)::get(null,"","PORT_652_COUNT",port_count[652]);
		     uvm_config_db #(int)::get(null,"","PORT_653_COUNT",port_count[653]);
		     uvm_config_db #(int)::get(null,"","PORT_654_COUNT",port_count[654]);
		     uvm_config_db #(int)::get(null,"","PORT_655_COUNT",port_count[655]);
		     uvm_config_db #(int)::get(null,"","PORT_656_COUNT",port_count[656]);
		     uvm_config_db #(int)::get(null,"","PORT_657_COUNT",port_count[657]);
		     uvm_config_db #(int)::get(null,"","PORT_658_COUNT",port_count[658]);
		     uvm_config_db #(int)::get(null,"","PORT_659_COUNT",port_count[659]);
		     uvm_config_db #(int)::get(null,"","PORT_660_COUNT",port_count[660]);
		     uvm_config_db #(int)::get(null,"","PORT_661_COUNT",port_count[661]);
		     uvm_config_db #(int)::get(null,"","PORT_662_COUNT",port_count[662]);
		     uvm_config_db #(int)::get(null,"","PORT_663_COUNT",port_count[663]);
		     uvm_config_db #(int)::get(null,"","PORT_664_COUNT",port_count[664]);
		     uvm_config_db #(int)::get(null,"","PORT_665_COUNT",port_count[665]);
		     uvm_config_db #(int)::get(null,"","PORT_666_COUNT",port_count[666]);
		     uvm_config_db #(int)::get(null,"","PORT_667_COUNT",port_count[667]);
		     uvm_config_db #(int)::get(null,"","PORT_668_COUNT",port_count[668]);
		     uvm_config_db #(int)::get(null,"","PORT_669_COUNT",port_count[669]);
		     uvm_config_db #(int)::get(null,"","PORT_670_COUNT",port_count[670]);
		     uvm_config_db #(int)::get(null,"","PORT_671_COUNT",port_count[671]);
		     uvm_config_db #(int)::get(null,"","PORT_672_COUNT",port_count[672]);
		     uvm_config_db #(int)::get(null,"","PORT_673_COUNT",port_count[673]);
		     uvm_config_db #(int)::get(null,"","PORT_674_COUNT",port_count[674]);
		     uvm_config_db #(int)::get(null,"","PORT_675_COUNT",port_count[675]);
		     uvm_config_db #(int)::get(null,"","PORT_676_COUNT",port_count[676]);
		     uvm_config_db #(int)::get(null,"","PORT_677_COUNT",port_count[677]);
		     uvm_config_db #(int)::get(null,"","PORT_678_COUNT",port_count[678]);
		     uvm_config_db #(int)::get(null,"","PORT_679_COUNT",port_count[679]);
		     uvm_config_db #(int)::get(null,"","PORT_680_COUNT",port_count[680]);
		     uvm_config_db #(int)::get(null,"","PORT_681_COUNT",port_count[681]);
		     uvm_config_db #(int)::get(null,"","PORT_682_COUNT",port_count[682]);
		     uvm_config_db #(int)::get(null,"","PORT_683_COUNT",port_count[683]);
		     uvm_config_db #(int)::get(null,"","PORT_684_COUNT",port_count[684]);
		     uvm_config_db #(int)::get(null,"","PORT_685_COUNT",port_count[685]);
		     uvm_config_db #(int)::get(null,"","PORT_686_COUNT",port_count[686]);
		     uvm_config_db #(int)::get(null,"","PORT_687_COUNT",port_count[687]);
		     uvm_config_db #(int)::get(null,"","PORT_688_COUNT",port_count[688]);
		     uvm_config_db #(int)::get(null,"","PORT_689_COUNT",port_count[689]);
		     uvm_config_db #(int)::get(null,"","PORT_690_COUNT",port_count[690]);
		     uvm_config_db #(int)::get(null,"","PORT_691_COUNT",port_count[691]);
		     uvm_config_db #(int)::get(null,"","PORT_692_COUNT",port_count[692]);
		     uvm_config_db #(int)::get(null,"","PORT_693_COUNT",port_count[693]);
		     uvm_config_db #(int)::get(null,"","PORT_694_COUNT",port_count[694]);
		     uvm_config_db #(int)::get(null,"","PORT_695_COUNT",port_count[695]);
		     uvm_config_db #(int)::get(null,"","PORT_696_COUNT",port_count[696]);
		     uvm_config_db #(int)::get(null,"","PORT_697_COUNT",port_count[697]);
		     uvm_config_db #(int)::get(null,"","PORT_698_COUNT",port_count[698]);
		     uvm_config_db #(int)::get(null,"","PORT_699_COUNT",port_count[699]);
		     uvm_config_db #(int)::get(null,"","PORT_700_COUNT",port_count[700]);
		     uvm_config_db #(int)::get(null,"","PORT_701_COUNT",port_count[701]);
		     uvm_config_db #(int)::get(null,"","PORT_702_COUNT",port_count[702]);
		     uvm_config_db #(int)::get(null,"","PORT_703_COUNT",port_count[703]);
		     uvm_config_db #(int)::get(null,"","PORT_704_COUNT",port_count[704]);
		     uvm_config_db #(int)::get(null,"","PORT_705_COUNT",port_count[705]);
		     uvm_config_db #(int)::get(null,"","PORT_706_COUNT",port_count[706]);
		     uvm_config_db #(int)::get(null,"","PORT_707_COUNT",port_count[707]);
		     uvm_config_db #(int)::get(null,"","PORT_708_COUNT",port_count[708]);
		     uvm_config_db #(int)::get(null,"","PORT_709_COUNT",port_count[709]);
		     uvm_config_db #(int)::get(null,"","PORT_710_COUNT",port_count[710]);
		     uvm_config_db #(int)::get(null,"","PORT_711_COUNT",port_count[711]);
		     uvm_config_db #(int)::get(null,"","PORT_712_COUNT",port_count[712]);
		     uvm_config_db #(int)::get(null,"","PORT_713_COUNT",port_count[713]);
		     uvm_config_db #(int)::get(null,"","PORT_714_COUNT",port_count[714]);
		     uvm_config_db #(int)::get(null,"","PORT_715_COUNT",port_count[715]);
		     uvm_config_db #(int)::get(null,"","PORT_716_COUNT",port_count[716]);
		     uvm_config_db #(int)::get(null,"","PORT_717_COUNT",port_count[717]);
		     uvm_config_db #(int)::get(null,"","PORT_718_COUNT",port_count[718]);
		     uvm_config_db #(int)::get(null,"","PORT_719_COUNT",port_count[719]);
		     uvm_config_db #(int)::get(null,"","PORT_720_COUNT",port_count[720]);
		     uvm_config_db #(int)::get(null,"","PORT_721_COUNT",port_count[721]);
		     uvm_config_db #(int)::get(null,"","PORT_722_COUNT",port_count[722]);
		     uvm_config_db #(int)::get(null,"","PORT_723_COUNT",port_count[723]);
		     uvm_config_db #(int)::get(null,"","PORT_724_COUNT",port_count[724]);
		     uvm_config_db #(int)::get(null,"","PORT_725_COUNT",port_count[725]);
		     uvm_config_db #(int)::get(null,"","PORT_726_COUNT",port_count[726]);
		     uvm_config_db #(int)::get(null,"","PORT_727_COUNT",port_count[727]);
		     uvm_config_db #(int)::get(null,"","PORT_728_COUNT",port_count[728]);
		     uvm_config_db #(int)::get(null,"","PORT_729_COUNT",port_count[729]);
		     uvm_config_db #(int)::get(null,"","PORT_730_COUNT",port_count[730]);
		     uvm_config_db #(int)::get(null,"","PORT_731_COUNT",port_count[731]);
		     uvm_config_db #(int)::get(null,"","PORT_732_COUNT",port_count[732]);
		     uvm_config_db #(int)::get(null,"","PORT_733_COUNT",port_count[733]);
		     uvm_config_db #(int)::get(null,"","PORT_734_COUNT",port_count[734]);
		     uvm_config_db #(int)::get(null,"","PORT_735_COUNT",port_count[735]);
		     uvm_config_db #(int)::get(null,"","PORT_736_COUNT",port_count[736]);
		     uvm_config_db #(int)::get(null,"","PORT_737_COUNT",port_count[737]);
		     uvm_config_db #(int)::get(null,"","PORT_738_COUNT",port_count[738]);
		     uvm_config_db #(int)::get(null,"","PORT_739_COUNT",port_count[739]);
		     uvm_config_db #(int)::get(null,"","PORT_740_COUNT",port_count[740]);
		     uvm_config_db #(int)::get(null,"","PORT_741_COUNT",port_count[741]);
		     uvm_config_db #(int)::get(null,"","PORT_742_COUNT",port_count[742]);
		     uvm_config_db #(int)::get(null,"","PORT_743_COUNT",port_count[743]);
		     uvm_config_db #(int)::get(null,"","PORT_744_COUNT",port_count[744]);
		     uvm_config_db #(int)::get(null,"","PORT_745_COUNT",port_count[745]);
		     uvm_config_db #(int)::get(null,"","PORT_746_COUNT",port_count[746]);
		     uvm_config_db #(int)::get(null,"","PORT_747_COUNT",port_count[747]);
		     uvm_config_db #(int)::get(null,"","PORT_748_COUNT",port_count[748]);
		     uvm_config_db #(int)::get(null,"","PORT_749_COUNT",port_count[749]);
		     uvm_config_db #(int)::get(null,"","PORT_750_COUNT",port_count[750]);
		     uvm_config_db #(int)::get(null,"","PORT_751_COUNT",port_count[751]);
		     uvm_config_db #(int)::get(null,"","PORT_752_COUNT",port_count[752]);
		     uvm_config_db #(int)::get(null,"","PORT_753_COUNT",port_count[753]);
		     uvm_config_db #(int)::get(null,"","PORT_754_COUNT",port_count[754]);
		     uvm_config_db #(int)::get(null,"","PORT_755_COUNT",port_count[755]);
		     uvm_config_db #(int)::get(null,"","PORT_756_COUNT",port_count[756]);
		     uvm_config_db #(int)::get(null,"","PORT_757_COUNT",port_count[757]);
		     uvm_config_db #(int)::get(null,"","PORT_758_COUNT",port_count[758]);
		     uvm_config_db #(int)::get(null,"","PORT_759_COUNT",port_count[759]);
		     uvm_config_db #(int)::get(null,"","PORT_760_COUNT",port_count[760]);
		     uvm_config_db #(int)::get(null,"","PORT_761_COUNT",port_count[761]);
		     uvm_config_db #(int)::get(null,"","PORT_762_COUNT",port_count[762]);
		     uvm_config_db #(int)::get(null,"","PORT_763_COUNT",port_count[763]);
		     uvm_config_db #(int)::get(null,"","PORT_764_COUNT",port_count[764]);
		     uvm_config_db #(int)::get(null,"","PORT_765_COUNT",port_count[765]);
		     uvm_config_db #(int)::get(null,"","PORT_766_COUNT",port_count[766]);
		     uvm_config_db #(int)::get(null,"","PORT_767_COUNT",port_count[767]);
		     uvm_config_db #(int)::get(null,"","PORT_768_COUNT",port_count[768]);
		     uvm_config_db #(int)::get(null,"","PORT_769_COUNT",port_count[769]);
		     uvm_config_db #(int)::get(null,"","PORT_770_COUNT",port_count[770]);
		     uvm_config_db #(int)::get(null,"","PORT_771_COUNT",port_count[771]);
		     uvm_config_db #(int)::get(null,"","PORT_772_COUNT",port_count[772]);
		     uvm_config_db #(int)::get(null,"","PORT_773_COUNT",port_count[773]);
		     uvm_config_db #(int)::get(null,"","PORT_774_COUNT",port_count[774]);
		     uvm_config_db #(int)::get(null,"","PORT_775_COUNT",port_count[775]);
		     uvm_config_db #(int)::get(null,"","PORT_776_COUNT",port_count[776]);
		     uvm_config_db #(int)::get(null,"","PORT_777_COUNT",port_count[777]);
		     uvm_config_db #(int)::get(null,"","PORT_778_COUNT",port_count[778]);
		     uvm_config_db #(int)::get(null,"","PORT_779_COUNT",port_count[779]);
		     uvm_config_db #(int)::get(null,"","PORT_780_COUNT",port_count[780]);
		     uvm_config_db #(int)::get(null,"","PORT_781_COUNT",port_count[781]);
		     uvm_config_db #(int)::get(null,"","PORT_782_COUNT",port_count[782]);
		     uvm_config_db #(int)::get(null,"","PORT_783_COUNT",port_count[783]);
		     uvm_config_db #(int)::get(null,"","PORT_784_COUNT",port_count[784]);
		     uvm_config_db #(int)::get(null,"","PORT_785_COUNT",port_count[785]);
		     uvm_config_db #(int)::get(null,"","PORT_786_COUNT",port_count[786]);
		     uvm_config_db #(int)::get(null,"","PORT_787_COUNT",port_count[787]);
		     uvm_config_db #(int)::get(null,"","PORT_788_COUNT",port_count[788]);
		     uvm_config_db #(int)::get(null,"","PORT_789_COUNT",port_count[789]);
		     uvm_config_db #(int)::get(null,"","PORT_790_COUNT",port_count[790]);
		     uvm_config_db #(int)::get(null,"","PORT_791_COUNT",port_count[791]);
		     uvm_config_db #(int)::get(null,"","PORT_792_COUNT",port_count[792]);
		     uvm_config_db #(int)::get(null,"","PORT_793_COUNT",port_count[793]);
		     uvm_config_db #(int)::get(null,"","PORT_794_COUNT",port_count[794]);
		     uvm_config_db #(int)::get(null,"","PORT_795_COUNT",port_count[795]);
		     uvm_config_db #(int)::get(null,"","PORT_796_COUNT",port_count[796]);
		     uvm_config_db #(int)::get(null,"","PORT_797_COUNT",port_count[797]);
		     uvm_config_db #(int)::get(null,"","PORT_798_COUNT",port_count[798]);
		     uvm_config_db #(int)::get(null,"","PORT_799_COUNT",port_count[799]);
		     uvm_config_db #(int)::get(null,"","PORT_800_COUNT",port_count[800]);
		     uvm_config_db #(int)::get(null,"","PORT_801_COUNT",port_count[801]);
		     uvm_config_db #(int)::get(null,"","PORT_802_COUNT",port_count[802]);
		     uvm_config_db #(int)::get(null,"","PORT_803_COUNT",port_count[803]);
		     uvm_config_db #(int)::get(null,"","PORT_804_COUNT",port_count[804]);
		     uvm_config_db #(int)::get(null,"","PORT_805_COUNT",port_count[805]);
		     uvm_config_db #(int)::get(null,"","PORT_806_COUNT",port_count[806]);
		     uvm_config_db #(int)::get(null,"","PORT_807_COUNT",port_count[807]);
		     uvm_config_db #(int)::get(null,"","PORT_808_COUNT",port_count[808]);
		     uvm_config_db #(int)::get(null,"","PORT_809_COUNT",port_count[809]);
		     uvm_config_db #(int)::get(null,"","PORT_810_COUNT",port_count[810]);
		     uvm_config_db #(int)::get(null,"","PORT_811_COUNT",port_count[811]);
		     uvm_config_db #(int)::get(null,"","PORT_812_COUNT",port_count[812]);
		     uvm_config_db #(int)::get(null,"","PORT_813_COUNT",port_count[813]);
		     uvm_config_db #(int)::get(null,"","PORT_814_COUNT",port_count[814]);
		     uvm_config_db #(int)::get(null,"","PORT_815_COUNT",port_count[815]);
		     uvm_config_db #(int)::get(null,"","PORT_816_COUNT",port_count[816]);
		     uvm_config_db #(int)::get(null,"","PORT_817_COUNT",port_count[817]);
		     uvm_config_db #(int)::get(null,"","PORT_818_COUNT",port_count[818]);
		     uvm_config_db #(int)::get(null,"","PORT_819_COUNT",port_count[819]);
		     uvm_config_db #(int)::get(null,"","PORT_820_COUNT",port_count[820]);
		     uvm_config_db #(int)::get(null,"","PORT_821_COUNT",port_count[821]);
		     uvm_config_db #(int)::get(null,"","PORT_822_COUNT",port_count[822]);
		     uvm_config_db #(int)::get(null,"","PORT_823_COUNT",port_count[823]);
		     uvm_config_db #(int)::get(null,"","PORT_824_COUNT",port_count[824]);
		     uvm_config_db #(int)::get(null,"","PORT_825_COUNT",port_count[825]);
		     uvm_config_db #(int)::get(null,"","PORT_826_COUNT",port_count[826]);
		     uvm_config_db #(int)::get(null,"","PORT_827_COUNT",port_count[827]);
		     uvm_config_db #(int)::get(null,"","PORT_828_COUNT",port_count[828]);
		     uvm_config_db #(int)::get(null,"","PORT_829_COUNT",port_count[829]);
		     uvm_config_db #(int)::get(null,"","PORT_830_COUNT",port_count[830]);
		     uvm_config_db #(int)::get(null,"","PORT_831_COUNT",port_count[831]);
		     uvm_config_db #(int)::get(null,"","PORT_832_COUNT",port_count[832]);
		     uvm_config_db #(int)::get(null,"","PORT_833_COUNT",port_count[833]);
		     uvm_config_db #(int)::get(null,"","PORT_834_COUNT",port_count[834]);
		     uvm_config_db #(int)::get(null,"","PORT_835_COUNT",port_count[835]);
		     uvm_config_db #(int)::get(null,"","PORT_836_COUNT",port_count[836]);
		     uvm_config_db #(int)::get(null,"","PORT_837_COUNT",port_count[837]);
		     uvm_config_db #(int)::get(null,"","PORT_838_COUNT",port_count[838]);
		     uvm_config_db #(int)::get(null,"","PORT_839_COUNT",port_count[839]);
		     uvm_config_db #(int)::get(null,"","PORT_840_COUNT",port_count[840]);
		     uvm_config_db #(int)::get(null,"","PORT_841_COUNT",port_count[841]);
		     uvm_config_db #(int)::get(null,"","PORT_842_COUNT",port_count[842]);
		     uvm_config_db #(int)::get(null,"","PORT_843_COUNT",port_count[843]);
		     uvm_config_db #(int)::get(null,"","PORT_844_COUNT",port_count[844]);
		     uvm_config_db #(int)::get(null,"","PORT_845_COUNT",port_count[845]);
		     uvm_config_db #(int)::get(null,"","PORT_846_COUNT",port_count[846]);
		     uvm_config_db #(int)::get(null,"","PORT_847_COUNT",port_count[847]);
		     uvm_config_db #(int)::get(null,"","PORT_848_COUNT",port_count[848]);
		     uvm_config_db #(int)::get(null,"","PORT_849_COUNT",port_count[849]);
		     uvm_config_db #(int)::get(null,"","PORT_850_COUNT",port_count[850]);
		     uvm_config_db #(int)::get(null,"","PORT_851_COUNT",port_count[851]);
		     uvm_config_db #(int)::get(null,"","PORT_852_COUNT",port_count[852]);
		     uvm_config_db #(int)::get(null,"","PORT_853_COUNT",port_count[853]);
		     uvm_config_db #(int)::get(null,"","PORT_854_COUNT",port_count[854]);
		     uvm_config_db #(int)::get(null,"","PORT_855_COUNT",port_count[855]);
		     uvm_config_db #(int)::get(null,"","PORT_856_COUNT",port_count[856]);
		     uvm_config_db #(int)::get(null,"","PORT_857_COUNT",port_count[857]);
		     uvm_config_db #(int)::get(null,"","PORT_858_COUNT",port_count[858]);
		     uvm_config_db #(int)::get(null,"","PORT_859_COUNT",port_count[859]);
		     uvm_config_db #(int)::get(null,"","PORT_860_COUNT",port_count[860]);
		     uvm_config_db #(int)::get(null,"","PORT_861_COUNT",port_count[861]);
		     uvm_config_db #(int)::get(null,"","PORT_862_COUNT",port_count[862]);
		     uvm_config_db #(int)::get(null,"","PORT_863_COUNT",port_count[863]);
		     uvm_config_db #(int)::get(null,"","PORT_864_COUNT",port_count[864]);
		     uvm_config_db #(int)::get(null,"","PORT_865_COUNT",port_count[865]);
		     uvm_config_db #(int)::get(null,"","PORT_866_COUNT",port_count[866]);
		     uvm_config_db #(int)::get(null,"","PORT_867_COUNT",port_count[867]);
		     uvm_config_db #(int)::get(null,"","PORT_868_COUNT",port_count[868]);
		     uvm_config_db #(int)::get(null,"","PORT_869_COUNT",port_count[869]);
		     uvm_config_db #(int)::get(null,"","PORT_870_COUNT",port_count[870]);
		     uvm_config_db #(int)::get(null,"","PORT_871_COUNT",port_count[871]);
		     uvm_config_db #(int)::get(null,"","PORT_872_COUNT",port_count[872]);
		     uvm_config_db #(int)::get(null,"","PORT_873_COUNT",port_count[873]);
		     uvm_config_db #(int)::get(null,"","PORT_874_COUNT",port_count[874]);
		     uvm_config_db #(int)::get(null,"","PORT_875_COUNT",port_count[875]);
		     uvm_config_db #(int)::get(null,"","PORT_876_COUNT",port_count[876]);
		     uvm_config_db #(int)::get(null,"","PORT_877_COUNT",port_count[877]);
		     uvm_config_db #(int)::get(null,"","PORT_878_COUNT",port_count[878]);
		     uvm_config_db #(int)::get(null,"","PORT_879_COUNT",port_count[879]);
		     uvm_config_db #(int)::get(null,"","PORT_880_COUNT",port_count[880]);
		     uvm_config_db #(int)::get(null,"","PORT_881_COUNT",port_count[881]);
		     uvm_config_db #(int)::get(null,"","PORT_882_COUNT",port_count[882]);
		     uvm_config_db #(int)::get(null,"","PORT_883_COUNT",port_count[883]);
		     uvm_config_db #(int)::get(null,"","PORT_884_COUNT",port_count[884]);
		     uvm_config_db #(int)::get(null,"","PORT_885_COUNT",port_count[885]);
		     uvm_config_db #(int)::get(null,"","PORT_886_COUNT",port_count[886]);
		     uvm_config_db #(int)::get(null,"","PORT_887_COUNT",port_count[887]);
		     uvm_config_db #(int)::get(null,"","PORT_888_COUNT",port_count[888]);
		     uvm_config_db #(int)::get(null,"","PORT_889_COUNT",port_count[889]);
		     uvm_config_db #(int)::get(null,"","PORT_890_COUNT",port_count[890]);
		     uvm_config_db #(int)::get(null,"","PORT_891_COUNT",port_count[891]);
		     uvm_config_db #(int)::get(null,"","PORT_892_COUNT",port_count[892]);
		     uvm_config_db #(int)::get(null,"","PORT_893_COUNT",port_count[893]);
		     uvm_config_db #(int)::get(null,"","PORT_894_COUNT",port_count[894]);
		     uvm_config_db #(int)::get(null,"","PORT_895_COUNT",port_count[895]);
		     uvm_config_db #(int)::get(null,"","PORT_896_COUNT",port_count[896]);
		     uvm_config_db #(int)::get(null,"","PORT_897_COUNT",port_count[897]);
		     uvm_config_db #(int)::get(null,"","PORT_898_COUNT",port_count[898]);
		     uvm_config_db #(int)::get(null,"","PORT_899_COUNT",port_count[899]);
		     uvm_config_db #(int)::get(null,"","PORT_900_COUNT",port_count[900]);
		     uvm_config_db #(int)::get(null,"","PORT_901_COUNT",port_count[901]);
		     uvm_config_db #(int)::get(null,"","PORT_902_COUNT",port_count[902]);
		     uvm_config_db #(int)::get(null,"","PORT_903_COUNT",port_count[903]);
		     uvm_config_db #(int)::get(null,"","PORT_904_COUNT",port_count[904]);
		     uvm_config_db #(int)::get(null,"","PORT_905_COUNT",port_count[905]);
		     uvm_config_db #(int)::get(null,"","PORT_906_COUNT",port_count[906]);
		     uvm_config_db #(int)::get(null,"","PORT_907_COUNT",port_count[907]);
		     uvm_config_db #(int)::get(null,"","PORT_908_COUNT",port_count[908]);
		     uvm_config_db #(int)::get(null,"","PORT_909_COUNT",port_count[909]);
		     uvm_config_db #(int)::get(null,"","PORT_910_COUNT",port_count[910]);
		     uvm_config_db #(int)::get(null,"","PORT_911_COUNT",port_count[911]);
		     uvm_config_db #(int)::get(null,"","PORT_912_COUNT",port_count[912]);
		     uvm_config_db #(int)::get(null,"","PORT_913_COUNT",port_count[913]);
		     uvm_config_db #(int)::get(null,"","PORT_914_COUNT",port_count[914]);
		     uvm_config_db #(int)::get(null,"","PORT_915_COUNT",port_count[915]);
		     uvm_config_db #(int)::get(null,"","PORT_916_COUNT",port_count[916]);
		     uvm_config_db #(int)::get(null,"","PORT_917_COUNT",port_count[917]);
		     uvm_config_db #(int)::get(null,"","PORT_918_COUNT",port_count[918]);
		     uvm_config_db #(int)::get(null,"","PORT_919_COUNT",port_count[919]);
		     uvm_config_db #(int)::get(null,"","PORT_920_COUNT",port_count[920]);
		     uvm_config_db #(int)::get(null,"","PORT_921_COUNT",port_count[921]);
		     uvm_config_db #(int)::get(null,"","PORT_922_COUNT",port_count[922]);
		     uvm_config_db #(int)::get(null,"","PORT_923_COUNT",port_count[923]);
		     uvm_config_db #(int)::get(null,"","PORT_924_COUNT",port_count[924]);
		     uvm_config_db #(int)::get(null,"","PORT_925_COUNT",port_count[925]);
		     uvm_config_db #(int)::get(null,"","PORT_926_COUNT",port_count[926]);
		     uvm_config_db #(int)::get(null,"","PORT_927_COUNT",port_count[927]);
		     uvm_config_db #(int)::get(null,"","PORT_928_COUNT",port_count[928]);
		     uvm_config_db #(int)::get(null,"","PORT_929_COUNT",port_count[929]);
		     uvm_config_db #(int)::get(null,"","PORT_930_COUNT",port_count[930]);
		     uvm_config_db #(int)::get(null,"","PORT_931_COUNT",port_count[931]);
		     uvm_config_db #(int)::get(null,"","PORT_932_COUNT",port_count[932]);
		     uvm_config_db #(int)::get(null,"","PORT_933_COUNT",port_count[933]);
		     uvm_config_db #(int)::get(null,"","PORT_934_COUNT",port_count[934]);
		     uvm_config_db #(int)::get(null,"","PORT_935_COUNT",port_count[935]);
		     uvm_config_db #(int)::get(null,"","PORT_936_COUNT",port_count[936]);
		     uvm_config_db #(int)::get(null,"","PORT_937_COUNT",port_count[937]);
		     uvm_config_db #(int)::get(null,"","PORT_938_COUNT",port_count[938]);
		     uvm_config_db #(int)::get(null,"","PORT_939_COUNT",port_count[939]);
		     uvm_config_db #(int)::get(null,"","PORT_940_COUNT",port_count[940]);
		     uvm_config_db #(int)::get(null,"","PORT_941_COUNT",port_count[941]);
		     uvm_config_db #(int)::get(null,"","PORT_942_COUNT",port_count[942]);
		     uvm_config_db #(int)::get(null,"","PORT_943_COUNT",port_count[943]);
		     uvm_config_db #(int)::get(null,"","PORT_944_COUNT",port_count[944]);
		     uvm_config_db #(int)::get(null,"","PORT_945_COUNT",port_count[945]);
		     uvm_config_db #(int)::get(null,"","PORT_946_COUNT",port_count[946]);
		     uvm_config_db #(int)::get(null,"","PORT_947_COUNT",port_count[947]);
		     uvm_config_db #(int)::get(null,"","PORT_948_COUNT",port_count[948]);
		     uvm_config_db #(int)::get(null,"","PORT_949_COUNT",port_count[949]);
		     uvm_config_db #(int)::get(null,"","PORT_950_COUNT",port_count[950]);
		     uvm_config_db #(int)::get(null,"","PORT_951_COUNT",port_count[951]);
		     uvm_config_db #(int)::get(null,"","PORT_952_COUNT",port_count[952]);
		     uvm_config_db #(int)::get(null,"","PORT_953_COUNT",port_count[953]);
		     uvm_config_db #(int)::get(null,"","PORT_954_COUNT",port_count[954]);
		     uvm_config_db #(int)::get(null,"","PORT_955_COUNT",port_count[955]);
		     uvm_config_db #(int)::get(null,"","PORT_956_COUNT",port_count[956]);
		     uvm_config_db #(int)::get(null,"","PORT_957_COUNT",port_count[957]);
		     uvm_config_db #(int)::get(null,"","PORT_958_COUNT",port_count[958]);
		     uvm_config_db #(int)::get(null,"","PORT_959_COUNT",port_count[959]);
		     uvm_config_db #(int)::get(null,"","PORT_960_COUNT",port_count[960]);
		     uvm_config_db #(int)::get(null,"","PORT_961_COUNT",port_count[961]);
		     uvm_config_db #(int)::get(null,"","PORT_962_COUNT",port_count[962]);
		     uvm_config_db #(int)::get(null,"","PORT_963_COUNT",port_count[963]);
		     uvm_config_db #(int)::get(null,"","PORT_964_COUNT",port_count[964]);
		     uvm_config_db #(int)::get(null,"","PORT_965_COUNT",port_count[965]);
		     uvm_config_db #(int)::get(null,"","PORT_966_COUNT",port_count[966]);
		     uvm_config_db #(int)::get(null,"","PORT_967_COUNT",port_count[967]);
		     uvm_config_db #(int)::get(null,"","PORT_968_COUNT",port_count[968]);
		     uvm_config_db #(int)::get(null,"","PORT_969_COUNT",port_count[969]);
		     uvm_config_db #(int)::get(null,"","PORT_970_COUNT",port_count[970]);
		     uvm_config_db #(int)::get(null,"","PORT_971_COUNT",port_count[971]);
		     uvm_config_db #(int)::get(null,"","PORT_972_COUNT",port_count[972]);
		     uvm_config_db #(int)::get(null,"","PORT_973_COUNT",port_count[973]);
		     uvm_config_db #(int)::get(null,"","PORT_974_COUNT",port_count[974]);
		     uvm_config_db #(int)::get(null,"","PORT_975_COUNT",port_count[975]);
		     uvm_config_db #(int)::get(null,"","PORT_976_COUNT",port_count[976]);
		     uvm_config_db #(int)::get(null,"","PORT_977_COUNT",port_count[977]);
		     uvm_config_db #(int)::get(null,"","PORT_978_COUNT",port_count[978]);
		     uvm_config_db #(int)::get(null,"","PORT_979_COUNT",port_count[979]);
		     uvm_config_db #(int)::get(null,"","PORT_980_COUNT",port_count[980]);
		     uvm_config_db #(int)::get(null,"","PORT_981_COUNT",port_count[981]);
		     uvm_config_db #(int)::get(null,"","PORT_982_COUNT",port_count[982]);
		     uvm_config_db #(int)::get(null,"","PORT_983_COUNT",port_count[983]);
		     uvm_config_db #(int)::get(null,"","PORT_984_COUNT",port_count[984]);
		     uvm_config_db #(int)::get(null,"","PORT_985_COUNT",port_count[985]);
		     uvm_config_db #(int)::get(null,"","PORT_986_COUNT",port_count[986]);
		     uvm_config_db #(int)::get(null,"","PORT_987_COUNT",port_count[987]);
		     uvm_config_db #(int)::get(null,"","PORT_988_COUNT",port_count[988]);
		     uvm_config_db #(int)::get(null,"","PORT_989_COUNT",port_count[989]);
		     uvm_config_db #(int)::get(null,"","PORT_990_COUNT",port_count[990]);
		     uvm_config_db #(int)::get(null,"","PORT_991_COUNT",port_count[991]);
		     uvm_config_db #(int)::get(null,"","PORT_992_COUNT",port_count[992]);
		     uvm_config_db #(int)::get(null,"","PORT_993_COUNT",port_count[993]);
		     uvm_config_db #(int)::get(null,"","PORT_994_COUNT",port_count[994]);
		     uvm_config_db #(int)::get(null,"","PORT_995_COUNT",port_count[995]);
		     uvm_config_db #(int)::get(null,"","PORT_996_COUNT",port_count[996]);
		     uvm_config_db #(int)::get(null,"","PORT_997_COUNT",port_count[997]);
		     uvm_config_db #(int)::get(null,"","PORT_998_COUNT",port_count[998]);
		     uvm_config_db #(int)::get(null,"","PORT_999_COUNT",port_count[999]);
		     uvm_config_db #(int)::get(null,"","PORT_1000_COUNT",port_count[1000]);
		     uvm_config_db #(int)::get(null,"","PORT_1001_COUNT",port_count[1001]);
		     uvm_config_db #(int)::get(null,"","PORT_1002_COUNT",port_count[1002]);
		     uvm_config_db #(int)::get(null,"","PORT_1003_COUNT",port_count[1003]);
		     uvm_config_db #(int)::get(null,"","PORT_1004_COUNT",port_count[1004]);
		     uvm_config_db #(int)::get(null,"","PORT_1005_COUNT",port_count[1005]);
		     uvm_config_db #(int)::get(null,"","PORT_1006_COUNT",port_count[1006]);
		     uvm_config_db #(int)::get(null,"","PORT_1007_COUNT",port_count[1007]);
		     uvm_config_db #(int)::get(null,"","PORT_1008_COUNT",port_count[1008]);
		     uvm_config_db #(int)::get(null,"","PORT_1009_COUNT",port_count[1009]);
		     uvm_config_db #(int)::get(null,"","PORT_1010_COUNT",port_count[1010]);
		     uvm_config_db #(int)::get(null,"","PORT_1011_COUNT",port_count[1011]);
		     uvm_config_db #(int)::get(null,"","PORT_1012_COUNT",port_count[1012]);
		     uvm_config_db #(int)::get(null,"","PORT_1013_COUNT",port_count[1013]);
		     uvm_config_db #(int)::get(null,"","PORT_1014_COUNT",port_count[1014]);
		     uvm_config_db #(int)::get(null,"","PORT_1015_COUNT",port_count[1015]);
		     uvm_config_db #(int)::get(null,"","PORT_1016_COUNT",port_count[1016]);
		     uvm_config_db #(int)::get(null,"","PORT_1017_COUNT",port_count[1017]);
		     uvm_config_db #(int)::get(null,"","PORT_1018_COUNT",port_count[1018]);
		     uvm_config_db #(int)::get(null,"","PORT_1019_COUNT",port_count[1019]);
		     uvm_config_db #(int)::get(null,"","PORT_1020_COUNT",port_count[1020]);
		     uvm_config_db #(int)::get(null,"","PORT_1021_COUNT",port_count[1021]);
		     uvm_config_db #(int)::get(null,"","PORT_1022_COUNT",port_count[1022]);
		     uvm_config_db #(int)::get(null,"","PORT_1023_COUNT",port_count[1023]);
		     uvm_config_db #(int)::get(null,"","PORT_1024_COUNT",port_count[1024]);
		     uvm_config_db #(int)::get(null,"","PORT_1025_COUNT",port_count[1025]);
		     uvm_config_db #(int)::get(null,"","PORT_1026_COUNT",port_count[1026]);
		     uvm_config_db #(int)::get(null,"","PORT_1027_COUNT",port_count[1027]);
		     uvm_config_db #(int)::get(null,"","PORT_1028_COUNT",port_count[1028]);
		     uvm_config_db #(int)::get(null,"","PORT_1029_COUNT",port_count[1029]);
		     uvm_config_db #(int)::get(null,"","PORT_1030_COUNT",port_count[1030]);
		     uvm_config_db #(int)::get(null,"","PORT_1031_COUNT",port_count[1031]);
		     uvm_config_db #(int)::get(null,"","PORT_1032_COUNT",port_count[1032]);
		     uvm_config_db #(int)::get(null,"","PORT_1033_COUNT",port_count[1033]);
		     uvm_config_db #(int)::get(null,"","PORT_1034_COUNT",port_count[1034]);
		     uvm_config_db #(int)::get(null,"","PORT_1035_COUNT",port_count[1035]);
		     uvm_config_db #(int)::get(null,"","PORT_1036_COUNT",port_count[1036]);
		     uvm_config_db #(int)::get(null,"","PORT_1037_COUNT",port_count[1037]);
		     uvm_config_db #(int)::get(null,"","PORT_1038_COUNT",port_count[1038]);
		     uvm_config_db #(int)::get(null,"","PORT_1039_COUNT",port_count[1039]);
		     uvm_config_db #(int)::get(null,"","PORT_1040_COUNT",port_count[1040]);
		     uvm_config_db #(int)::get(null,"","PORT_1041_COUNT",port_count[1041]);
		     uvm_config_db #(int)::get(null,"","PORT_1042_COUNT",port_count[1042]);
		     uvm_config_db #(int)::get(null,"","PORT_1043_COUNT",port_count[1043]);
		     uvm_config_db #(int)::get(null,"","PORT_1044_COUNT",port_count[1044]);
		     uvm_config_db #(int)::get(null,"","PORT_1045_COUNT",port_count[1045]);
		     uvm_config_db #(int)::get(null,"","PORT_1046_COUNT",port_count[1046]);
		     uvm_config_db #(int)::get(null,"","PORT_1047_COUNT",port_count[1047]);
		     uvm_config_db #(int)::get(null,"","PORT_1048_COUNT",port_count[1048]);
		     uvm_config_db #(int)::get(null,"","PORT_1049_COUNT",port_count[1049]);
		     uvm_config_db #(int)::get(null,"","PORT_1050_COUNT",port_count[1050]);
		     uvm_config_db #(int)::get(null,"","PORT_1051_COUNT",port_count[1051]);
		     uvm_config_db #(int)::get(null,"","PORT_1052_COUNT",port_count[1052]);
		     uvm_config_db #(int)::get(null,"","PORT_1053_COUNT",port_count[1053]);
		     uvm_config_db #(int)::get(null,"","PORT_1054_COUNT",port_count[1054]);
		     uvm_config_db #(int)::get(null,"","PORT_1055_COUNT",port_count[1055]);
		     uvm_config_db #(int)::get(null,"","PORT_1056_COUNT",port_count[1056]);
		     uvm_config_db #(int)::get(null,"","PORT_1057_COUNT",port_count[1057]);
		     uvm_config_db #(int)::get(null,"","PORT_1058_COUNT",port_count[1058]);
		     uvm_config_db #(int)::get(null,"","PORT_1059_COUNT",port_count[1059]);
		     uvm_config_db #(int)::get(null,"","PORT_1060_COUNT",port_count[1060]);
		     uvm_config_db #(int)::get(null,"","PORT_1061_COUNT",port_count[1061]);
		     uvm_config_db #(int)::get(null,"","PORT_1062_COUNT",port_count[1062]);
		     uvm_config_db #(int)::get(null,"","PORT_1063_COUNT",port_count[1063]);
		     uvm_config_db #(int)::get(null,"","PORT_1064_COUNT",port_count[1064]);
		     uvm_config_db #(int)::get(null,"","PORT_1065_COUNT",port_count[1065]);
		     uvm_config_db #(int)::get(null,"","PORT_1066_COUNT",port_count[1066]);
		     uvm_config_db #(int)::get(null,"","PORT_1067_COUNT",port_count[1067]);
		     uvm_config_db #(int)::get(null,"","PORT_1068_COUNT",port_count[1068]);
		     uvm_config_db #(int)::get(null,"","PORT_1069_COUNT",port_count[1069]);
		     uvm_config_db #(int)::get(null,"","PORT_1070_COUNT",port_count[1070]);
		     uvm_config_db #(int)::get(null,"","PORT_1071_COUNT",port_count[1071]);
		     uvm_config_db #(int)::get(null,"","PORT_1072_COUNT",port_count[1072]);
		     uvm_config_db #(int)::get(null,"","PORT_1073_COUNT",port_count[1073]);
		     uvm_config_db #(int)::get(null,"","PORT_1074_COUNT",port_count[1074]);
		     uvm_config_db #(int)::get(null,"","PORT_1075_COUNT",port_count[1075]);
		     uvm_config_db #(int)::get(null,"","PORT_1076_COUNT",port_count[1076]);
		     uvm_config_db #(int)::get(null,"","PORT_1077_COUNT",port_count[1077]);
		     uvm_config_db #(int)::get(null,"","PORT_1078_COUNT",port_count[1078]);
		     uvm_config_db #(int)::get(null,"","PORT_1079_COUNT",port_count[1079]);
		     uvm_config_db #(int)::get(null,"","PORT_1080_COUNT",port_count[1080]);
		     uvm_config_db #(int)::get(null,"","PORT_1081_COUNT",port_count[1081]);
		     uvm_config_db #(int)::get(null,"","PORT_1082_COUNT",port_count[1082]);
		     uvm_config_db #(int)::get(null,"","PORT_1083_COUNT",port_count[1083]);
		     uvm_config_db #(int)::get(null,"","PORT_1084_COUNT",port_count[1084]);
		     uvm_config_db #(int)::get(null,"","PORT_1085_COUNT",port_count[1085]);
		     uvm_config_db #(int)::get(null,"","PORT_1086_COUNT",port_count[1086]);
		     uvm_config_db #(int)::get(null,"","PORT_1087_COUNT",port_count[1087]);
		     uvm_config_db #(int)::get(null,"","PORT_1088_COUNT",port_count[1088]);
		     uvm_config_db #(int)::get(null,"","PORT_1089_COUNT",port_count[1089]);
		     uvm_config_db #(int)::get(null,"","PORT_1090_COUNT",port_count[1090]);
		     uvm_config_db #(int)::get(null,"","PORT_1091_COUNT",port_count[1091]);
		     uvm_config_db #(int)::get(null,"","PORT_1092_COUNT",port_count[1092]);
		     uvm_config_db #(int)::get(null,"","PORT_1093_COUNT",port_count[1093]);
		     uvm_config_db #(int)::get(null,"","PORT_1094_COUNT",port_count[1094]);
		     uvm_config_db #(int)::get(null,"","PORT_1095_COUNT",port_count[1095]);
		     uvm_config_db #(int)::get(null,"","PORT_1096_COUNT",port_count[1096]);
		     uvm_config_db #(int)::get(null,"","PORT_1097_COUNT",port_count[1097]);
		     uvm_config_db #(int)::get(null,"","PORT_1098_COUNT",port_count[1098]);
		     uvm_config_db #(int)::get(null,"","PORT_1099_COUNT",port_count[1099]);
		     uvm_config_db #(int)::get(null,"","PORT_1100_COUNT",port_count[1100]);
		     uvm_config_db #(int)::get(null,"","PORT_1101_COUNT",port_count[1101]);
		     uvm_config_db #(int)::get(null,"","PORT_1102_COUNT",port_count[1102]);
		     uvm_config_db #(int)::get(null,"","PORT_1103_COUNT",port_count[1103]);
		     uvm_config_db #(int)::get(null,"","PORT_1104_COUNT",port_count[1104]);
		     uvm_config_db #(int)::get(null,"","PORT_1105_COUNT",port_count[1105]);
		     uvm_config_db #(int)::get(null,"","PORT_1106_COUNT",port_count[1106]);
		     uvm_config_db #(int)::get(null,"","PORT_1107_COUNT",port_count[1107]);
		     uvm_config_db #(int)::get(null,"","PORT_1108_COUNT",port_count[1108]);
		     uvm_config_db #(int)::get(null,"","PORT_1109_COUNT",port_count[1109]);
		     uvm_config_db #(int)::get(null,"","PORT_1110_COUNT",port_count[1110]);
		     uvm_config_db #(int)::get(null,"","PORT_1111_COUNT",port_count[1111]);
		     uvm_config_db #(int)::get(null,"","PORT_1112_COUNT",port_count[1112]);
		     uvm_config_db #(int)::get(null,"","PORT_1113_COUNT",port_count[1113]);
		     uvm_config_db #(int)::get(null,"","PORT_1114_COUNT",port_count[1114]);
		     uvm_config_db #(int)::get(null,"","PORT_1115_COUNT",port_count[1115]);
		     uvm_config_db #(int)::get(null,"","PORT_1116_COUNT",port_count[1116]);
		     uvm_config_db #(int)::get(null,"","PORT_1117_COUNT",port_count[1117]);
		     uvm_config_db #(int)::get(null,"","PORT_1118_COUNT",port_count[1118]);
		     uvm_config_db #(int)::get(null,"","PORT_1119_COUNT",port_count[1119]);
		     uvm_config_db #(int)::get(null,"","PORT_1120_COUNT",port_count[1120]);
		     uvm_config_db #(int)::get(null,"","PORT_1121_COUNT",port_count[1121]);
		     uvm_config_db #(int)::get(null,"","PORT_1122_COUNT",port_count[1122]);
		     uvm_config_db #(int)::get(null,"","PORT_1123_COUNT",port_count[1123]);
		     uvm_config_db #(int)::get(null,"","PORT_1124_COUNT",port_count[1124]);
		     uvm_config_db #(int)::get(null,"","PORT_1125_COUNT",port_count[1125]);
		     uvm_config_db #(int)::get(null,"","PORT_1126_COUNT",port_count[1126]);
		     uvm_config_db #(int)::get(null,"","PORT_1127_COUNT",port_count[1127]);
		     uvm_config_db #(int)::get(null,"","PORT_1128_COUNT",port_count[1128]);
		     uvm_config_db #(int)::get(null,"","PORT_1129_COUNT",port_count[1129]);
		     uvm_config_db #(int)::get(null,"","PORT_1130_COUNT",port_count[1130]);
		     uvm_config_db #(int)::get(null,"","PORT_1131_COUNT",port_count[1131]);
		     uvm_config_db #(int)::get(null,"","PORT_1132_COUNT",port_count[1132]);
		     uvm_config_db #(int)::get(null,"","PORT_1133_COUNT",port_count[1133]);
		     uvm_config_db #(int)::get(null,"","PORT_1134_COUNT",port_count[1134]);
		     uvm_config_db #(int)::get(null,"","PORT_1135_COUNT",port_count[1135]);
		     uvm_config_db #(int)::get(null,"","PORT_1136_COUNT",port_count[1136]);
		     uvm_config_db #(int)::get(null,"","PORT_1137_COUNT",port_count[1137]);
		     uvm_config_db #(int)::get(null,"","PORT_1138_COUNT",port_count[1138]);
		     uvm_config_db #(int)::get(null,"","PORT_1139_COUNT",port_count[1139]);
		     uvm_config_db #(int)::get(null,"","PORT_1140_COUNT",port_count[1140]);
		     uvm_config_db #(int)::get(null,"","PORT_1141_COUNT",port_count[1141]);
		     uvm_config_db #(int)::get(null,"","PORT_1142_COUNT",port_count[1142]);
		     uvm_config_db #(int)::get(null,"","PORT_1143_COUNT",port_count[1143]);
		     uvm_config_db #(int)::get(null,"","PORT_1144_COUNT",port_count[1144]);
		     uvm_config_db #(int)::get(null,"","PORT_1145_COUNT",port_count[1145]);
		     uvm_config_db #(int)::get(null,"","PORT_1146_COUNT",port_count[1146]);
		     uvm_config_db #(int)::get(null,"","PORT_1147_COUNT",port_count[1147]);
		     uvm_config_db #(int)::get(null,"","PORT_1148_COUNT",port_count[1148]);
		     uvm_config_db #(int)::get(null,"","PORT_1149_COUNT",port_count[1149]);
		     uvm_config_db #(int)::get(null,"","PORT_1150_COUNT",port_count[1150]);
		     uvm_config_db #(int)::get(null,"","PORT_1151_COUNT",port_count[1151]);
		     uvm_config_db #(int)::get(null,"","PORT_1152_COUNT",port_count[1152]);
		     uvm_config_db #(int)::get(null,"","PORT_1153_COUNT",port_count[1153]);
		     uvm_config_db #(int)::get(null,"","PORT_1154_COUNT",port_count[1154]);
		     uvm_config_db #(int)::get(null,"","PORT_1155_COUNT",port_count[1155]);
		     uvm_config_db #(int)::get(null,"","PORT_1156_COUNT",port_count[1156]);
		     uvm_config_db #(int)::get(null,"","PORT_1157_COUNT",port_count[1157]);
		     uvm_config_db #(int)::get(null,"","PORT_1158_COUNT",port_count[1158]);
		     uvm_config_db #(int)::get(null,"","PORT_1159_COUNT",port_count[1159]);
		     uvm_config_db #(int)::get(null,"","PORT_1160_COUNT",port_count[1160]);
		     uvm_config_db #(int)::get(null,"","PORT_1161_COUNT",port_count[1161]);
		     uvm_config_db #(int)::get(null,"","PORT_1162_COUNT",port_count[1162]);
		     uvm_config_db #(int)::get(null,"","PORT_1163_COUNT",port_count[1163]);
		     uvm_config_db #(int)::get(null,"","PORT_1164_COUNT",port_count[1164]);
		     uvm_config_db #(int)::get(null,"","PORT_1165_COUNT",port_count[1165]);
		     uvm_config_db #(int)::get(null,"","PORT_1166_COUNT",port_count[1166]);
		     uvm_config_db #(int)::get(null,"","PORT_1167_COUNT",port_count[1167]);
		     uvm_config_db #(int)::get(null,"","PORT_1168_COUNT",port_count[1168]);
		     uvm_config_db #(int)::get(null,"","PORT_1169_COUNT",port_count[1169]);
		     uvm_config_db #(int)::get(null,"","PORT_1170_COUNT",port_count[1170]);
		     uvm_config_db #(int)::get(null,"","PORT_1171_COUNT",port_count[1171]);
		     uvm_config_db #(int)::get(null,"","PORT_1172_COUNT",port_count[1172]);
		     uvm_config_db #(int)::get(null,"","PORT_1173_COUNT",port_count[1173]);
		     uvm_config_db #(int)::get(null,"","PORT_1174_COUNT",port_count[1174]);
		     uvm_config_db #(int)::get(null,"","PORT_1175_COUNT",port_count[1175]);
		     uvm_config_db #(int)::get(null,"","PORT_1176_COUNT",port_count[1176]);
		     uvm_config_db #(int)::get(null,"","PORT_1177_COUNT",port_count[1177]);
		     uvm_config_db #(int)::get(null,"","PORT_1178_COUNT",port_count[1178]);
		     uvm_config_db #(int)::get(null,"","PORT_1179_COUNT",port_count[1179]);
		     uvm_config_db #(int)::get(null,"","PORT_1180_COUNT",port_count[1180]);
		     uvm_config_db #(int)::get(null,"","PORT_1181_COUNT",port_count[1181]);
		     uvm_config_db #(int)::get(null,"","PORT_1182_COUNT",port_count[1182]);
		     uvm_config_db #(int)::get(null,"","PORT_1183_COUNT",port_count[1183]);
		     uvm_config_db #(int)::get(null,"","PORT_1184_COUNT",port_count[1184]);
		     uvm_config_db #(int)::get(null,"","PORT_1185_COUNT",port_count[1185]);
		     uvm_config_db #(int)::get(null,"","PORT_1186_COUNT",port_count[1186]);
		     uvm_config_db #(int)::get(null,"","PORT_1187_COUNT",port_count[1187]);
		     uvm_config_db #(int)::get(null,"","PORT_1188_COUNT",port_count[1188]);
		     uvm_config_db #(int)::get(null,"","PORT_1189_COUNT",port_count[1189]);
		     uvm_config_db #(int)::get(null,"","PORT_1190_COUNT",port_count[1190]);
		     uvm_config_db #(int)::get(null,"","PORT_1191_COUNT",port_count[1191]);
		     uvm_config_db #(int)::get(null,"","PORT_1192_COUNT",port_count[1192]);
		     uvm_config_db #(int)::get(null,"","PORT_1193_COUNT",port_count[1193]);
		     uvm_config_db #(int)::get(null,"","PORT_1194_COUNT",port_count[1194]);
		     uvm_config_db #(int)::get(null,"","PORT_1195_COUNT",port_count[1195]);
		     uvm_config_db #(int)::get(null,"","PORT_1196_COUNT",port_count[1196]);
		     uvm_config_db #(int)::get(null,"","PORT_1197_COUNT",port_count[1197]);
		     uvm_config_db #(int)::get(null,"","PORT_1198_COUNT",port_count[1198]);
		     uvm_config_db #(int)::get(null,"","PORT_1199_COUNT",port_count[1199]);
		     uvm_config_db #(int)::get(null,"","PORT_1200_COUNT",port_count[1200]);
		     uvm_config_db #(int)::get(null,"","PORT_1201_COUNT",port_count[1201]);
		     uvm_config_db #(int)::get(null,"","PORT_1202_COUNT",port_count[1202]);
		     uvm_config_db #(int)::get(null,"","PORT_1203_COUNT",port_count[1203]);
		     uvm_config_db #(int)::get(null,"","PORT_1204_COUNT",port_count[1204]);
		     uvm_config_db #(int)::get(null,"","PORT_1205_COUNT",port_count[1205]);
		     uvm_config_db #(int)::get(null,"","PORT_1206_COUNT",port_count[1206]);
		     uvm_config_db #(int)::get(null,"","PORT_1207_COUNT",port_count[1207]);
		     uvm_config_db #(int)::get(null,"","PORT_1208_COUNT",port_count[1208]);
		     uvm_config_db #(int)::get(null,"","PORT_1209_COUNT",port_count[1209]);
		     uvm_config_db #(int)::get(null,"","PORT_1210_COUNT",port_count[1210]);
		     uvm_config_db #(int)::get(null,"","PORT_1211_COUNT",port_count[1211]);
		     uvm_config_db #(int)::get(null,"","PORT_1212_COUNT",port_count[1212]);
		     uvm_config_db #(int)::get(null,"","PORT_1213_COUNT",port_count[1213]);
		     uvm_config_db #(int)::get(null,"","PORT_1214_COUNT",port_count[1214]);
		     uvm_config_db #(int)::get(null,"","PORT_1215_COUNT",port_count[1215]);
		     uvm_config_db #(int)::get(null,"","PORT_1216_COUNT",port_count[1216]);
		     uvm_config_db #(int)::get(null,"","PORT_1217_COUNT",port_count[1217]);
		     uvm_config_db #(int)::get(null,"","PORT_1218_COUNT",port_count[1218]);
		     uvm_config_db #(int)::get(null,"","PORT_1219_COUNT",port_count[1219]);
		     uvm_config_db #(int)::get(null,"","PORT_1220_COUNT",port_count[1220]);
		     uvm_config_db #(int)::get(null,"","PORT_1221_COUNT",port_count[1221]);
		     uvm_config_db #(int)::get(null,"","PORT_1222_COUNT",port_count[1222]);
		     uvm_config_db #(int)::get(null,"","PORT_1223_COUNT",port_count[1223]);
		     uvm_config_db #(int)::get(null,"","PORT_1224_COUNT",port_count[1224]);
		     uvm_config_db #(int)::get(null,"","PORT_1225_COUNT",port_count[1225]);
		     uvm_config_db #(int)::get(null,"","PORT_1226_COUNT",port_count[1226]);
		     uvm_config_db #(int)::get(null,"","PORT_1227_COUNT",port_count[1227]);
		     uvm_config_db #(int)::get(null,"","PORT_1228_COUNT",port_count[1228]);
		     uvm_config_db #(int)::get(null,"","PORT_1229_COUNT",port_count[1229]);
		     uvm_config_db #(int)::get(null,"","PORT_1230_COUNT",port_count[1230]);
		     uvm_config_db #(int)::get(null,"","PORT_1231_COUNT",port_count[1231]);
		     uvm_config_db #(int)::get(null,"","PORT_1232_COUNT",port_count[1232]);
		     uvm_config_db #(int)::get(null,"","PORT_1233_COUNT",port_count[1233]);
		     uvm_config_db #(int)::get(null,"","PORT_1234_COUNT",port_count[1234]);
		     uvm_config_db #(int)::get(null,"","PORT_1235_COUNT",port_count[1235]);
		     uvm_config_db #(int)::get(null,"","PORT_1236_COUNT",port_count[1236]);
		     uvm_config_db #(int)::get(null,"","PORT_1237_COUNT",port_count[1237]);
		     uvm_config_db #(int)::get(null,"","PORT_1238_COUNT",port_count[1238]);
		     uvm_config_db #(int)::get(null,"","PORT_1239_COUNT",port_count[1239]);
		     uvm_config_db #(int)::get(null,"","PORT_1240_COUNT",port_count[1240]);
		     uvm_config_db #(int)::get(null,"","PORT_1241_COUNT",port_count[1241]);
		     uvm_config_db #(int)::get(null,"","PORT_1242_COUNT",port_count[1242]);
		     uvm_config_db #(int)::get(null,"","PORT_1243_COUNT",port_count[1243]);
		     uvm_config_db #(int)::get(null,"","PORT_1244_COUNT",port_count[1244]);
		     uvm_config_db #(int)::get(null,"","PORT_1245_COUNT",port_count[1245]);
		     uvm_config_db #(int)::get(null,"","PORT_1246_COUNT",port_count[1246]);
		     uvm_config_db #(int)::get(null,"","PORT_1247_COUNT",port_count[1247]);
		     uvm_config_db #(int)::get(null,"","PORT_1248_COUNT",port_count[1248]);
		     uvm_config_db #(int)::get(null,"","PORT_1249_COUNT",port_count[1249]);
		     uvm_config_db #(int)::get(null,"","PORT_1250_COUNT",port_count[1250]);
		     uvm_config_db #(int)::get(null,"","PORT_1251_COUNT",port_count[1251]);
		     uvm_config_db #(int)::get(null,"","PORT_1252_COUNT",port_count[1252]);
		     uvm_config_db #(int)::get(null,"","PORT_1253_COUNT",port_count[1253]);
		     uvm_config_db #(int)::get(null,"","PORT_1254_COUNT",port_count[1254]);
		     uvm_config_db #(int)::get(null,"","PORT_1255_COUNT",port_count[1255]);
		     uvm_config_db #(int)::get(null,"","PORT_1256_COUNT",port_count[1256]);
		     uvm_config_db #(int)::get(null,"","PORT_1257_COUNT",port_count[1257]);
		     uvm_config_db #(int)::get(null,"","PORT_1258_COUNT",port_count[1258]);
		     uvm_config_db #(int)::get(null,"","PORT_1259_COUNT",port_count[1259]);
		     uvm_config_db #(int)::get(null,"","PORT_1260_COUNT",port_count[1260]);
		     uvm_config_db #(int)::get(null,"","PORT_1261_COUNT",port_count[1261]);
		     uvm_config_db #(int)::get(null,"","PORT_1262_COUNT",port_count[1262]);
		     uvm_config_db #(int)::get(null,"","PORT_1263_COUNT",port_count[1263]);
		     uvm_config_db #(int)::get(null,"","PORT_1264_COUNT",port_count[1264]);
		     uvm_config_db #(int)::get(null,"","PORT_1265_COUNT",port_count[1265]);
		     uvm_config_db #(int)::get(null,"","PORT_1266_COUNT",port_count[1266]);
		     uvm_config_db #(int)::get(null,"","PORT_1267_COUNT",port_count[1267]);
		     uvm_config_db #(int)::get(null,"","PORT_1268_COUNT",port_count[1268]);
		     uvm_config_db #(int)::get(null,"","PORT_1269_COUNT",port_count[1269]);
		     uvm_config_db #(int)::get(null,"","PORT_1270_COUNT",port_count[1270]);
		     uvm_config_db #(int)::get(null,"","PORT_1271_COUNT",port_count[1271]);
		     uvm_config_db #(int)::get(null,"","PORT_1272_COUNT",port_count[1272]);
		     uvm_config_db #(int)::get(null,"","PORT_1273_COUNT",port_count[1273]);
		     uvm_config_db #(int)::get(null,"","PORT_1274_COUNT",port_count[1274]);
		     uvm_config_db #(int)::get(null,"","PORT_1275_COUNT",port_count[1275]);
		     uvm_config_db #(int)::get(null,"","PORT_1276_COUNT",port_count[1276]);
		     uvm_config_db #(int)::get(null,"","PORT_1277_COUNT",port_count[1277]);
		     uvm_config_db #(int)::get(null,"","PORT_1278_COUNT",port_count[1278]);
		     uvm_config_db #(int)::get(null,"","PORT_1279_COUNT",port_count[1279]);
		     uvm_config_db #(int)::get(null,"","PORT_1280_COUNT",port_count[1280]);
		     uvm_config_db #(int)::get(null,"","PORT_1281_COUNT",port_count[1281]);
		     uvm_config_db #(int)::get(null,"","PORT_1282_COUNT",port_count[1282]);
		     uvm_config_db #(int)::get(null,"","PORT_1283_COUNT",port_count[1283]);
		     uvm_config_db #(int)::get(null,"","PORT_1284_COUNT",port_count[1284]);
		     uvm_config_db #(int)::get(null,"","PORT_1285_COUNT",port_count[1285]);
		     uvm_config_db #(int)::get(null,"","PORT_1286_COUNT",port_count[1286]);
		     uvm_config_db #(int)::get(null,"","PORT_1287_COUNT",port_count[1287]);
		     uvm_config_db #(int)::get(null,"","PORT_1288_COUNT",port_count[1288]);
		     uvm_config_db #(int)::get(null,"","PORT_1289_COUNT",port_count[1289]);
		     uvm_config_db #(int)::get(null,"","PORT_1290_COUNT",port_count[1290]);
		     uvm_config_db #(int)::get(null,"","PORT_1291_COUNT",port_count[1291]);
		     uvm_config_db #(int)::get(null,"","PORT_1292_COUNT",port_count[1292]);
		     uvm_config_db #(int)::get(null,"","PORT_1293_COUNT",port_count[1293]);
		     uvm_config_db #(int)::get(null,"","PORT_1294_COUNT",port_count[1294]);
		     uvm_config_db #(int)::get(null,"","PORT_1295_COUNT",port_count[1295]);
		     uvm_config_db #(int)::get(null,"","PORT_1296_COUNT",port_count[1296]);
		     uvm_config_db #(int)::get(null,"","PORT_1297_COUNT",port_count[1297]);
		     uvm_config_db #(int)::get(null,"","PORT_1298_COUNT",port_count[1298]);
		     uvm_config_db #(int)::get(null,"","PORT_1299_COUNT",port_count[1299]);
		     uvm_config_db #(int)::get(null,"","PORT_1300_COUNT",port_count[1300]);
		     uvm_config_db #(int)::get(null,"","PORT_1301_COUNT",port_count[1301]);
		     uvm_config_db #(int)::get(null,"","PORT_1302_COUNT",port_count[1302]);
		     uvm_config_db #(int)::get(null,"","PORT_1303_COUNT",port_count[1303]);
		     uvm_config_db #(int)::get(null,"","PORT_1304_COUNT",port_count[1304]);
		     uvm_config_db #(int)::get(null,"","PORT_1305_COUNT",port_count[1305]);
		     uvm_config_db #(int)::get(null,"","PORT_1306_COUNT",port_count[1306]);
		     uvm_config_db #(int)::get(null,"","PORT_1307_COUNT",port_count[1307]);
		     uvm_config_db #(int)::get(null,"","PORT_1308_COUNT",port_count[1308]);
		     uvm_config_db #(int)::get(null,"","PORT_1309_COUNT",port_count[1309]);
		     uvm_config_db #(int)::get(null,"","PORT_1310_COUNT",port_count[1310]);
		     uvm_config_db #(int)::get(null,"","PORT_1311_COUNT",port_count[1311]);
		     uvm_config_db #(int)::get(null,"","PORT_1312_COUNT",port_count[1312]);
		     uvm_config_db #(int)::get(null,"","PORT_1313_COUNT",port_count[1313]);
		     uvm_config_db #(int)::get(null,"","PORT_1314_COUNT",port_count[1314]);
		     uvm_config_db #(int)::get(null,"","PORT_1315_COUNT",port_count[1315]);
		     uvm_config_db #(int)::get(null,"","PORT_1316_COUNT",port_count[1316]);
		     uvm_config_db #(int)::get(null,"","PORT_1317_COUNT",port_count[1317]);
		     uvm_config_db #(int)::get(null,"","PORT_1318_COUNT",port_count[1318]);
		     uvm_config_db #(int)::get(null,"","PORT_1319_COUNT",port_count[1319]);
		     uvm_config_db #(int)::get(null,"","PORT_1320_COUNT",port_count[1320]);
		     uvm_config_db #(int)::get(null,"","PORT_1321_COUNT",port_count[1321]);
		     uvm_config_db #(int)::get(null,"","PORT_1322_COUNT",port_count[1322]);
		     uvm_config_db #(int)::get(null,"","PORT_1323_COUNT",port_count[1323]);
		     uvm_config_db #(int)::get(null,"","PORT_1324_COUNT",port_count[1324]);
		     uvm_config_db #(int)::get(null,"","PORT_1325_COUNT",port_count[1325]);
		     uvm_config_db #(int)::get(null,"","PORT_1326_COUNT",port_count[1326]);
		     uvm_config_db #(int)::get(null,"","PORT_1327_COUNT",port_count[1327]);
		     uvm_config_db #(int)::get(null,"","PORT_1328_COUNT",port_count[1328]);
		     uvm_config_db #(int)::get(null,"","PORT_1329_COUNT",port_count[1329]);
		     uvm_config_db #(int)::get(null,"","PORT_1330_COUNT",port_count[1330]);
		     uvm_config_db #(int)::get(null,"","PORT_1331_COUNT",port_count[1331]);
		     uvm_config_db #(int)::get(null,"","PORT_1332_COUNT",port_count[1332]);
		     uvm_config_db #(int)::get(null,"","PORT_1333_COUNT",port_count[1333]);
		     uvm_config_db #(int)::get(null,"","PORT_1334_COUNT",port_count[1334]);
		     uvm_config_db #(int)::get(null,"","PORT_1335_COUNT",port_count[1335]);
		     uvm_config_db #(int)::get(null,"","PORT_1336_COUNT",port_count[1336]);
		     uvm_config_db #(int)::get(null,"","PORT_1337_COUNT",port_count[1337]);
		     uvm_config_db #(int)::get(null,"","PORT_1338_COUNT",port_count[1338]);
		     uvm_config_db #(int)::get(null,"","PORT_1339_COUNT",port_count[1339]);
		     uvm_config_db #(int)::get(null,"","PORT_1340_COUNT",port_count[1340]);
		     uvm_config_db #(int)::get(null,"","PORT_1341_COUNT",port_count[1341]);
		     uvm_config_db #(int)::get(null,"","PORT_1342_COUNT",port_count[1342]);
		     uvm_config_db #(int)::get(null,"","PORT_1343_COUNT",port_count[1343]);
		     uvm_config_db #(int)::get(null,"","PORT_1344_COUNT",port_count[1344]);
		     uvm_config_db #(int)::get(null,"","PORT_1345_COUNT",port_count[1345]);
		     uvm_config_db #(int)::get(null,"","PORT_1346_COUNT",port_count[1346]);
		     uvm_config_db #(int)::get(null,"","PORT_1347_COUNT",port_count[1347]);
		     uvm_config_db #(int)::get(null,"","PORT_1348_COUNT",port_count[1348]);
		     uvm_config_db #(int)::get(null,"","PORT_1349_COUNT",port_count[1349]);
		     uvm_config_db #(int)::get(null,"","PORT_1350_COUNT",port_count[1350]);
		     uvm_config_db #(int)::get(null,"","PORT_1351_COUNT",port_count[1351]);
		     uvm_config_db #(int)::get(null,"","PORT_1352_COUNT",port_count[1352]);
		     uvm_config_db #(int)::get(null,"","PORT_1353_COUNT",port_count[1353]);
		     uvm_config_db #(int)::get(null,"","PORT_1354_COUNT",port_count[1354]);
		     uvm_config_db #(int)::get(null,"","PORT_1355_COUNT",port_count[1355]);
		     uvm_config_db #(int)::get(null,"","PORT_1356_COUNT",port_count[1356]);
		     uvm_config_db #(int)::get(null,"","PORT_1357_COUNT",port_count[1357]);
		     uvm_config_db #(int)::get(null,"","PORT_1358_COUNT",port_count[1358]);
		     uvm_config_db #(int)::get(null,"","PORT_1359_COUNT",port_count[1359]);
		     uvm_config_db #(int)::get(null,"","PORT_1360_COUNT",port_count[1360]);
		     uvm_config_db #(int)::get(null,"","PORT_1361_COUNT",port_count[1361]);
		     uvm_config_db #(int)::get(null,"","PORT_1362_COUNT",port_count[1362]);
		     uvm_config_db #(int)::get(null,"","PORT_1363_COUNT",port_count[1363]);
		     uvm_config_db #(int)::get(null,"","PORT_1364_COUNT",port_count[1364]);
		     uvm_config_db #(int)::get(null,"","PORT_1365_COUNT",port_count[1365]);
		     uvm_config_db #(int)::get(null,"","PORT_1366_COUNT",port_count[1366]);
		     uvm_config_db #(int)::get(null,"","PORT_1367_COUNT",port_count[1367]);
		     uvm_config_db #(int)::get(null,"","PORT_1368_COUNT",port_count[1368]);
		     uvm_config_db #(int)::get(null,"","PORT_1369_COUNT",port_count[1369]);
		     uvm_config_db #(int)::get(null,"","PORT_1370_COUNT",port_count[1370]);
		     uvm_config_db #(int)::get(null,"","PORT_1371_COUNT",port_count[1371]);
		     uvm_config_db #(int)::get(null,"","PORT_1372_COUNT",port_count[1372]);
		     uvm_config_db #(int)::get(null,"","PORT_1373_COUNT",port_count[1373]);
		     uvm_config_db #(int)::get(null,"","PORT_1374_COUNT",port_count[1374]);
		     uvm_config_db #(int)::get(null,"","PORT_1375_COUNT",port_count[1375]);
		     uvm_config_db #(int)::get(null,"","PORT_1376_COUNT",port_count[1376]);
		     uvm_config_db #(int)::get(null,"","PORT_1377_COUNT",port_count[1377]);
		     uvm_config_db #(int)::get(null,"","PORT_1378_COUNT",port_count[1378]);
		     uvm_config_db #(int)::get(null,"","PORT_1379_COUNT",port_count[1379]);
		     uvm_config_db #(int)::get(null,"","PORT_1380_COUNT",port_count[1380]);
		     uvm_config_db #(int)::get(null,"","PORT_1381_COUNT",port_count[1381]);
		     uvm_config_db #(int)::get(null,"","PORT_1382_COUNT",port_count[1382]);
		     uvm_config_db #(int)::get(null,"","PORT_1383_COUNT",port_count[1383]);
		     uvm_config_db #(int)::get(null,"","PORT_1384_COUNT",port_count[1384]);
		     uvm_config_db #(int)::get(null,"","PORT_1385_COUNT",port_count[1385]);
		     uvm_config_db #(int)::get(null,"","PORT_1386_COUNT",port_count[1386]);
		     uvm_config_db #(int)::get(null,"","PORT_1387_COUNT",port_count[1387]);
		     uvm_config_db #(int)::get(null,"","PORT_1388_COUNT",port_count[1388]);
		     uvm_config_db #(int)::get(null,"","PORT_1389_COUNT",port_count[1389]);
		     uvm_config_db #(int)::get(null,"","PORT_1390_COUNT",port_count[1390]);
		     uvm_config_db #(int)::get(null,"","PORT_1391_COUNT",port_count[1391]);
		     uvm_config_db #(int)::get(null,"","PORT_1392_COUNT",port_count[1392]);
		     uvm_config_db #(int)::get(null,"","PORT_1393_COUNT",port_count[1393]);
		     uvm_config_db #(int)::get(null,"","PORT_1394_COUNT",port_count[1394]);
		     uvm_config_db #(int)::get(null,"","PORT_1395_COUNT",port_count[1395]);
		     uvm_config_db #(int)::get(null,"","PORT_1396_COUNT",port_count[1396]);
		     uvm_config_db #(int)::get(null,"","PORT_1397_COUNT",port_count[1397]);
		     uvm_config_db #(int)::get(null,"","PORT_1398_COUNT",port_count[1398]);
		     uvm_config_db #(int)::get(null,"","PORT_1399_COUNT",port_count[1399]);
		     uvm_config_db #(int)::get(null,"","PORT_1400_COUNT",port_count[1400]);
		     uvm_config_db #(int)::get(null,"","PORT_1401_COUNT",port_count[1401]);
		     uvm_config_db #(int)::get(null,"","PORT_1402_COUNT",port_count[1402]);
		     uvm_config_db #(int)::get(null,"","PORT_1403_COUNT",port_count[1403]);
		     uvm_config_db #(int)::get(null,"","PORT_1404_COUNT",port_count[1404]);
		     uvm_config_db #(int)::get(null,"","PORT_1405_COUNT",port_count[1405]);
		     uvm_config_db #(int)::get(null,"","PORT_1406_COUNT",port_count[1406]);
		     uvm_config_db #(int)::get(null,"","PORT_1407_COUNT",port_count[1407]);
		     uvm_config_db #(int)::get(null,"","PORT_1408_COUNT",port_count[1408]);
		     uvm_config_db #(int)::get(null,"","PORT_1409_COUNT",port_count[1409]);
		     uvm_config_db #(int)::get(null,"","PORT_1410_COUNT",port_count[1410]);
		     uvm_config_db #(int)::get(null,"","PORT_1411_COUNT",port_count[1411]);
		     uvm_config_db #(int)::get(null,"","PORT_1412_COUNT",port_count[1412]);
		     uvm_config_db #(int)::get(null,"","PORT_1413_COUNT",port_count[1413]);
		     uvm_config_db #(int)::get(null,"","PORT_1414_COUNT",port_count[1414]);
		     uvm_config_db #(int)::get(null,"","PORT_1415_COUNT",port_count[1415]);
		     uvm_config_db #(int)::get(null,"","PORT_1416_COUNT",port_count[1416]);
		     uvm_config_db #(int)::get(null,"","PORT_1417_COUNT",port_count[1417]);
		     uvm_config_db #(int)::get(null,"","PORT_1418_COUNT",port_count[1418]);
		     uvm_config_db #(int)::get(null,"","PORT_1419_COUNT",port_count[1419]);
		     uvm_config_db #(int)::get(null,"","PORT_1420_COUNT",port_count[1420]);
		     uvm_config_db #(int)::get(null,"","PORT_1421_COUNT",port_count[1421]);
		     uvm_config_db #(int)::get(null,"","PORT_1422_COUNT",port_count[1422]);
		     uvm_config_db #(int)::get(null,"","PORT_1423_COUNT",port_count[1423]);
		     uvm_config_db #(int)::get(null,"","PORT_1424_COUNT",port_count[1424]);
		     uvm_config_db #(int)::get(null,"","PORT_1425_COUNT",port_count[1425]);
		     uvm_config_db #(int)::get(null,"","PORT_1426_COUNT",port_count[1426]);
		     uvm_config_db #(int)::get(null,"","PORT_1427_COUNT",port_count[1427]);
		     uvm_config_db #(int)::get(null,"","PORT_1428_COUNT",port_count[1428]);
		     uvm_config_db #(int)::get(null,"","PORT_1429_COUNT",port_count[1429]);
		     uvm_config_db #(int)::get(null,"","PORT_1430_COUNT",port_count[1430]);
		     uvm_config_db #(int)::get(null,"","PORT_1431_COUNT",port_count[1431]);
		     uvm_config_db #(int)::get(null,"","PORT_1432_COUNT",port_count[1432]);
		     uvm_config_db #(int)::get(null,"","PORT_1433_COUNT",port_count[1433]);
		     uvm_config_db #(int)::get(null,"","PORT_1434_COUNT",port_count[1434]);
		     uvm_config_db #(int)::get(null,"","PORT_1435_COUNT",port_count[1435]);
		     uvm_config_db #(int)::get(null,"","PORT_1436_COUNT",port_count[1436]);
		     uvm_config_db #(int)::get(null,"","PORT_1437_COUNT",port_count[1437]);
		     uvm_config_db #(int)::get(null,"","PORT_1438_COUNT",port_count[1438]);
		     uvm_config_db #(int)::get(null,"","PORT_1439_COUNT",port_count[1439]);
		     uvm_config_db #(int)::get(null,"","PORT_1440_COUNT",port_count[1440]);
		     uvm_config_db #(int)::get(null,"","PORT_1441_COUNT",port_count[1441]);
		     uvm_config_db #(int)::get(null,"","PORT_1442_COUNT",port_count[1442]);
		     uvm_config_db #(int)::get(null,"","PORT_1443_COUNT",port_count[1443]);
		     uvm_config_db #(int)::get(null,"","PORT_1444_COUNT",port_count[1444]);
		     uvm_config_db #(int)::get(null,"","PORT_1445_COUNT",port_count[1445]);
		     uvm_config_db #(int)::get(null,"","PORT_1446_COUNT",port_count[1446]);
		     uvm_config_db #(int)::get(null,"","PORT_1447_COUNT",port_count[1447]);
		     uvm_config_db #(int)::get(null,"","PORT_1448_COUNT",port_count[1448]);
		     uvm_config_db #(int)::get(null,"","PORT_1449_COUNT",port_count[1449]);
		     uvm_config_db #(int)::get(null,"","PORT_1450_COUNT",port_count[1450]);
		     uvm_config_db #(int)::get(null,"","PORT_1451_COUNT",port_count[1451]);
		     uvm_config_db #(int)::get(null,"","PORT_1452_COUNT",port_count[1452]);
		     uvm_config_db #(int)::get(null,"","PORT_1453_COUNT",port_count[1453]);
		     uvm_config_db #(int)::get(null,"","PORT_1454_COUNT",port_count[1454]);
		     uvm_config_db #(int)::get(null,"","PORT_1455_COUNT",port_count[1455]);
		     uvm_config_db #(int)::get(null,"","PORT_1456_COUNT",port_count[1456]);
		     uvm_config_db #(int)::get(null,"","PORT_1457_COUNT",port_count[1457]);
		     uvm_config_db #(int)::get(null,"","PORT_1458_COUNT",port_count[1458]);
		     uvm_config_db #(int)::get(null,"","PORT_1459_COUNT",port_count[1459]);
		     uvm_config_db #(int)::get(null,"","PORT_1460_COUNT",port_count[1460]);
		     uvm_config_db #(int)::get(null,"","PORT_1461_COUNT",port_count[1461]);
		     uvm_config_db #(int)::get(null,"","PORT_1462_COUNT",port_count[1462]);
		     uvm_config_db #(int)::get(null,"","PORT_1463_COUNT",port_count[1463]);
		     uvm_config_db #(int)::get(null,"","PORT_1464_COUNT",port_count[1464]);
		     uvm_config_db #(int)::get(null,"","PORT_1465_COUNT",port_count[1465]);
		     uvm_config_db #(int)::get(null,"","PORT_1466_COUNT",port_count[1466]);
		     uvm_config_db #(int)::get(null,"","PORT_1467_COUNT",port_count[1467]);
		     uvm_config_db #(int)::get(null,"","PORT_1468_COUNT",port_count[1468]);
		     uvm_config_db #(int)::get(null,"","PORT_1469_COUNT",port_count[1469]);
		     uvm_config_db #(int)::get(null,"","PORT_1470_COUNT",port_count[1470]);
		     uvm_config_db #(int)::get(null,"","PORT_1471_COUNT",port_count[1471]);
		     uvm_config_db #(int)::get(null,"","PORT_1472_COUNT",port_count[1472]);
		     uvm_config_db #(int)::get(null,"","PORT_1473_COUNT",port_count[1473]);
		     uvm_config_db #(int)::get(null,"","PORT_1474_COUNT",port_count[1474]);
		     uvm_config_db #(int)::get(null,"","PORT_1475_COUNT",port_count[1475]);
		     uvm_config_db #(int)::get(null,"","PORT_1476_COUNT",port_count[1476]);
		     uvm_config_db #(int)::get(null,"","PORT_1477_COUNT",port_count[1477]);
		     uvm_config_db #(int)::get(null,"","PORT_1478_COUNT",port_count[1478]);
		     uvm_config_db #(int)::get(null,"","PORT_1479_COUNT",port_count[1479]);
		     uvm_config_db #(int)::get(null,"","PORT_1480_COUNT",port_count[1480]);
		     uvm_config_db #(int)::get(null,"","PORT_1481_COUNT",port_count[1481]);
		     uvm_config_db #(int)::get(null,"","PORT_1482_COUNT",port_count[1482]);
		     uvm_config_db #(int)::get(null,"","PORT_1483_COUNT",port_count[1483]);
		     uvm_config_db #(int)::get(null,"","PORT_1484_COUNT",port_count[1484]);
		     uvm_config_db #(int)::get(null,"","PORT_1485_COUNT",port_count[1485]);
		     uvm_config_db #(int)::get(null,"","PORT_1486_COUNT",port_count[1486]);
		     uvm_config_db #(int)::get(null,"","PORT_1487_COUNT",port_count[1487]);
		     uvm_config_db #(int)::get(null,"","PORT_1488_COUNT",port_count[1488]);
		     uvm_config_db #(int)::get(null,"","PORT_1489_COUNT",port_count[1489]);
		     uvm_config_db #(int)::get(null,"","PORT_1490_COUNT",port_count[1490]);
		     uvm_config_db #(int)::get(null,"","PORT_1491_COUNT",port_count[1491]);
		     uvm_config_db #(int)::get(null,"","PORT_1492_COUNT",port_count[1492]);
		     uvm_config_db #(int)::get(null,"","PORT_1493_COUNT",port_count[1493]);
		     uvm_config_db #(int)::get(null,"","PORT_1494_COUNT",port_count[1494]);
		     uvm_config_db #(int)::get(null,"","PORT_1495_COUNT",port_count[1495]);
		     uvm_config_db #(int)::get(null,"","PORT_1496_COUNT",port_count[1496]);
		     uvm_config_db #(int)::get(null,"","PORT_1497_COUNT",port_count[1497]);
		     uvm_config_db #(int)::get(null,"","PORT_1498_COUNT",port_count[1498]);
		     uvm_config_db #(int)::get(null,"","PORT_1499_COUNT",port_count[1499]);
		     uvm_config_db #(int)::get(null,"","PORT_1500_COUNT",port_count[1500]);
		     uvm_config_db #(int)::get(null,"","PORT_1501_COUNT",port_count[1501]);
		     uvm_config_db #(int)::get(null,"","PORT_1502_COUNT",port_count[1502]);
		     uvm_config_db #(int)::get(null,"","PORT_1503_COUNT",port_count[1503]);
		     uvm_config_db #(int)::get(null,"","PORT_1504_COUNT",port_count[1504]);
		     uvm_config_db #(int)::get(null,"","PORT_1505_COUNT",port_count[1505]);
		     uvm_config_db #(int)::get(null,"","PORT_1506_COUNT",port_count[1506]);
		     uvm_config_db #(int)::get(null,"","PORT_1507_COUNT",port_count[1507]);
		     uvm_config_db #(int)::get(null,"","PORT_1508_COUNT",port_count[1508]);
		     uvm_config_db #(int)::get(null,"","PORT_1509_COUNT",port_count[1509]);
		     uvm_config_db #(int)::get(null,"","PORT_1510_COUNT",port_count[1510]);
		     uvm_config_db #(int)::get(null,"","PORT_1511_COUNT",port_count[1511]);
		     uvm_config_db #(int)::get(null,"","PORT_1512_COUNT",port_count[1512]);
		     uvm_config_db #(int)::get(null,"","PORT_1513_COUNT",port_count[1513]);
		     uvm_config_db #(int)::get(null,"","PORT_1514_COUNT",port_count[1514]);
		     uvm_config_db #(int)::get(null,"","PORT_1515_COUNT",port_count[1515]);
		     uvm_config_db #(int)::get(null,"","PORT_1516_COUNT",port_count[1516]);
		     uvm_config_db #(int)::get(null,"","PORT_1517_COUNT",port_count[1517]);
		     uvm_config_db #(int)::get(null,"","PORT_1518_COUNT",port_count[1518]);
		     uvm_config_db #(int)::get(null,"","PORT_1519_COUNT",port_count[1519]);
		     uvm_config_db #(int)::get(null,"","PORT_1520_COUNT",port_count[1520]);
		     uvm_config_db #(int)::get(null,"","PORT_1521_COUNT",port_count[1521]);
		     uvm_config_db #(int)::get(null,"","PORT_1522_COUNT",port_count[1522]);
		     uvm_config_db #(int)::get(null,"","PORT_1523_COUNT",port_count[1523]);
		     uvm_config_db #(int)::get(null,"","PORT_1524_COUNT",port_count[1524]);
		     uvm_config_db #(int)::get(null,"","PORT_1525_COUNT",port_count[1525]);
		     uvm_config_db #(int)::get(null,"","PORT_1526_COUNT",port_count[1526]);
		     uvm_config_db #(int)::get(null,"","PORT_1527_COUNT",port_count[1527]);
		     uvm_config_db #(int)::get(null,"","PORT_1528_COUNT",port_count[1528]);
		     uvm_config_db #(int)::get(null,"","PORT_1529_COUNT",port_count[1529]);
		     uvm_config_db #(int)::get(null,"","PORT_1530_COUNT",port_count[1530]);
		     uvm_config_db #(int)::get(null,"","PORT_1531_COUNT",port_count[1531]);
		     uvm_config_db #(int)::get(null,"","PORT_1532_COUNT",port_count[1532]);
		     uvm_config_db #(int)::get(null,"","PORT_1533_COUNT",port_count[1533]);
		     uvm_config_db #(int)::get(null,"","PORT_1534_COUNT",port_count[1534]);
		     uvm_config_db #(int)::get(null,"","PORT_1535_COUNT",port_count[1535]);
		     uvm_config_db #(int)::get(null,"","PORT_1536_COUNT",port_count[1536]);
		     uvm_config_db #(int)::get(null,"","PORT_1537_COUNT",port_count[1537]);
		     uvm_config_db #(int)::get(null,"","PORT_1538_COUNT",port_count[1538]);
		     uvm_config_db #(int)::get(null,"","PORT_1539_COUNT",port_count[1539]);
		     uvm_config_db #(int)::get(null,"","PORT_1540_COUNT",port_count[1540]);
		     uvm_config_db #(int)::get(null,"","PORT_1541_COUNT",port_count[1541]);
		     uvm_config_db #(int)::get(null,"","PORT_1542_COUNT",port_count[1542]);
		     uvm_config_db #(int)::get(null,"","PORT_1543_COUNT",port_count[1543]);
		     uvm_config_db #(int)::get(null,"","PORT_1544_COUNT",port_count[1544]);
		     uvm_config_db #(int)::get(null,"","PORT_1545_COUNT",port_count[1545]);
		     uvm_config_db #(int)::get(null,"","PORT_1546_COUNT",port_count[1546]);
		     uvm_config_db #(int)::get(null,"","PORT_1547_COUNT",port_count[1547]);
		     uvm_config_db #(int)::get(null,"","PORT_1548_COUNT",port_count[1548]);
		     uvm_config_db #(int)::get(null,"","PORT_1549_COUNT",port_count[1549]);
		     uvm_config_db #(int)::get(null,"","PORT_1550_COUNT",port_count[1550]);
		     uvm_config_db #(int)::get(null,"","PORT_1551_COUNT",port_count[1551]);
		     uvm_config_db #(int)::get(null,"","PORT_1552_COUNT",port_count[1552]);
		     uvm_config_db #(int)::get(null,"","PORT_1553_COUNT",port_count[1553]);
		     uvm_config_db #(int)::get(null,"","PORT_1554_COUNT",port_count[1554]);
		     uvm_config_db #(int)::get(null,"","PORT_1555_COUNT",port_count[1555]);
		     uvm_config_db #(int)::get(null,"","PORT_1556_COUNT",port_count[1556]);
		     uvm_config_db #(int)::get(null,"","PORT_1557_COUNT",port_count[1557]);
		     uvm_config_db #(int)::get(null,"","PORT_1558_COUNT",port_count[1558]);
		     uvm_config_db #(int)::get(null,"","PORT_1559_COUNT",port_count[1559]);
		     uvm_config_db #(int)::get(null,"","PORT_1560_COUNT",port_count[1560]);
		     uvm_config_db #(int)::get(null,"","PORT_1561_COUNT",port_count[1561]);
		     uvm_config_db #(int)::get(null,"","PORT_1562_COUNT",port_count[1562]);
		     uvm_config_db #(int)::get(null,"","PORT_1563_COUNT",port_count[1563]);
		     uvm_config_db #(int)::get(null,"","PORT_1564_COUNT",port_count[1564]);
		     uvm_config_db #(int)::get(null,"","PORT_1565_COUNT",port_count[1565]);
		     uvm_config_db #(int)::get(null,"","PORT_1566_COUNT",port_count[1566]);
		     uvm_config_db #(int)::get(null,"","PORT_1567_COUNT",port_count[1567]);
		     uvm_config_db #(int)::get(null,"","PORT_1568_COUNT",port_count[1568]);
		     uvm_config_db #(int)::get(null,"","PORT_1569_COUNT",port_count[1569]);
		     uvm_config_db #(int)::get(null,"","PORT_1570_COUNT",port_count[1570]);
		     uvm_config_db #(int)::get(null,"","PORT_1571_COUNT",port_count[1571]);
		     uvm_config_db #(int)::get(null,"","PORT_1572_COUNT",port_count[1572]);
		     uvm_config_db #(int)::get(null,"","PORT_1573_COUNT",port_count[1573]);
		     uvm_config_db #(int)::get(null,"","PORT_1574_COUNT",port_count[1574]);
		     uvm_config_db #(int)::get(null,"","PORT_1575_COUNT",port_count[1575]);
		     uvm_config_db #(int)::get(null,"","PORT_1576_COUNT",port_count[1576]);
		     uvm_config_db #(int)::get(null,"","PORT_1577_COUNT",port_count[1577]);
		     uvm_config_db #(int)::get(null,"","PORT_1578_COUNT",port_count[1578]);
		     uvm_config_db #(int)::get(null,"","PORT_1579_COUNT",port_count[1579]);
		     uvm_config_db #(int)::get(null,"","PORT_1580_COUNT",port_count[1580]);
		     uvm_config_db #(int)::get(null,"","PORT_1581_COUNT",port_count[1581]);
		     uvm_config_db #(int)::get(null,"","PORT_1582_COUNT",port_count[1582]);
		     uvm_config_db #(int)::get(null,"","PORT_1583_COUNT",port_count[1583]);
		     uvm_config_db #(int)::get(null,"","PORT_1584_COUNT",port_count[1584]);
		     uvm_config_db #(int)::get(null,"","PORT_1585_COUNT",port_count[1585]);
		     uvm_config_db #(int)::get(null,"","PORT_1586_COUNT",port_count[1586]);
		     uvm_config_db #(int)::get(null,"","PORT_1587_COUNT",port_count[1587]);
		     uvm_config_db #(int)::get(null,"","PORT_1588_COUNT",port_count[1588]);
		     uvm_config_db #(int)::get(null,"","PORT_1589_COUNT",port_count[1589]);
		     uvm_config_db #(int)::get(null,"","PORT_1590_COUNT",port_count[1590]);
		     uvm_config_db #(int)::get(null,"","PORT_1591_COUNT",port_count[1591]);
		     uvm_config_db #(int)::get(null,"","PORT_1592_COUNT",port_count[1592]);
		     uvm_config_db #(int)::get(null,"","PORT_1593_COUNT",port_count[1593]);
		     uvm_config_db #(int)::get(null,"","PORT_1594_COUNT",port_count[1594]);
		     uvm_config_db #(int)::get(null,"","PORT_1595_COUNT",port_count[1595]);
		     uvm_config_db #(int)::get(null,"","PORT_1596_COUNT",port_count[1596]);
		     uvm_config_db #(int)::get(null,"","PORT_1597_COUNT",port_count[1597]);
		     uvm_config_db #(int)::get(null,"","PORT_1598_COUNT",port_count[1598]);
		     uvm_config_db #(int)::get(null,"","PORT_1599_COUNT",port_count[1599]);
		     uvm_config_db #(int)::get(null,"","PORT_1600_COUNT",port_count[1600]);
		     uvm_config_db #(int)::get(null,"","PORT_1601_COUNT",port_count[1601]);
		     uvm_config_db #(int)::get(null,"","PORT_1602_COUNT",port_count[1602]);
		     uvm_config_db #(int)::get(null,"","PORT_1603_COUNT",port_count[1603]);
		     uvm_config_db #(int)::get(null,"","PORT_1604_COUNT",port_count[1604]);
		     uvm_config_db #(int)::get(null,"","PORT_1605_COUNT",port_count[1605]);
		     uvm_config_db #(int)::get(null,"","PORT_1606_COUNT",port_count[1606]);
		     uvm_config_db #(int)::get(null,"","PORT_1607_COUNT",port_count[1607]);
		     uvm_config_db #(int)::get(null,"","PORT_1608_COUNT",port_count[1608]);
		     uvm_config_db #(int)::get(null,"","PORT_1609_COUNT",port_count[1609]);
		     uvm_config_db #(int)::get(null,"","PORT_1610_COUNT",port_count[1610]);
		     uvm_config_db #(int)::get(null,"","PORT_1611_COUNT",port_count[1611]);
		     uvm_config_db #(int)::get(null,"","PORT_1612_COUNT",port_count[1612]);
		     uvm_config_db #(int)::get(null,"","PORT_1613_COUNT",port_count[1613]);
		     uvm_config_db #(int)::get(null,"","PORT_1614_COUNT",port_count[1614]);
		     uvm_config_db #(int)::get(null,"","PORT_1615_COUNT",port_count[1615]);
		     uvm_config_db #(int)::get(null,"","PORT_1616_COUNT",port_count[1616]);
		     uvm_config_db #(int)::get(null,"","PORT_1617_COUNT",port_count[1617]);
		     uvm_config_db #(int)::get(null,"","PORT_1618_COUNT",port_count[1618]);
		     uvm_config_db #(int)::get(null,"","PORT_1619_COUNT",port_count[1619]);
		     uvm_config_db #(int)::get(null,"","PORT_1620_COUNT",port_count[1620]);
		     uvm_config_db #(int)::get(null,"","PORT_1621_COUNT",port_count[1621]);
		     uvm_config_db #(int)::get(null,"","PORT_1622_COUNT",port_count[1622]);
		     uvm_config_db #(int)::get(null,"","PORT_1623_COUNT",port_count[1623]);
		     uvm_config_db #(int)::get(null,"","PORT_1624_COUNT",port_count[1624]);
		     uvm_config_db #(int)::get(null,"","PORT_1625_COUNT",port_count[1625]);
		     uvm_config_db #(int)::get(null,"","PORT_1626_COUNT",port_count[1626]);
		     uvm_config_db #(int)::get(null,"","PORT_1627_COUNT",port_count[1627]);
		     uvm_config_db #(int)::get(null,"","PORT_1628_COUNT",port_count[1628]);
		     uvm_config_db #(int)::get(null,"","PORT_1629_COUNT",port_count[1629]);
		     uvm_config_db #(int)::get(null,"","PORT_1630_COUNT",port_count[1630]);
		     uvm_config_db #(int)::get(null,"","PORT_1631_COUNT",port_count[1631]);
		     uvm_config_db #(int)::get(null,"","PORT_1632_COUNT",port_count[1632]);
		     uvm_config_db #(int)::get(null,"","PORT_1633_COUNT",port_count[1633]);
		     uvm_config_db #(int)::get(null,"","PORT_1634_COUNT",port_count[1634]);
		     uvm_config_db #(int)::get(null,"","PORT_1635_COUNT",port_count[1635]);
		     uvm_config_db #(int)::get(null,"","PORT_1636_COUNT",port_count[1636]);
		     uvm_config_db #(int)::get(null,"","PORT_1637_COUNT",port_count[1637]);
		     uvm_config_db #(int)::get(null,"","PORT_1638_COUNT",port_count[1638]);
		     uvm_config_db #(int)::get(null,"","PORT_1639_COUNT",port_count[1639]);
		     uvm_config_db #(int)::get(null,"","PORT_1640_COUNT",port_count[1640]);
		     uvm_config_db #(int)::get(null,"","PORT_1641_COUNT",port_count[1641]);
		     uvm_config_db #(int)::get(null,"","PORT_1642_COUNT",port_count[1642]);
		     uvm_config_db #(int)::get(null,"","PORT_1643_COUNT",port_count[1643]);
		     uvm_config_db #(int)::get(null,"","PORT_1644_COUNT",port_count[1644]);
		     uvm_config_db #(int)::get(null,"","PORT_1645_COUNT",port_count[1645]);
		     uvm_config_db #(int)::get(null,"","PORT_1646_COUNT",port_count[1646]);
		     uvm_config_db #(int)::get(null,"","PORT_1647_COUNT",port_count[1647]);
		     uvm_config_db #(int)::get(null,"","PORT_1648_COUNT",port_count[1648]);
		     uvm_config_db #(int)::get(null,"","PORT_1649_COUNT",port_count[1649]);
		     uvm_config_db #(int)::get(null,"","PORT_1650_COUNT",port_count[1650]);
		     uvm_config_db #(int)::get(null,"","PORT_1651_COUNT",port_count[1651]);
		     uvm_config_db #(int)::get(null,"","PORT_1652_COUNT",port_count[1652]);
		     uvm_config_db #(int)::get(null,"","PORT_1653_COUNT",port_count[1653]);
		     uvm_config_db #(int)::get(null,"","PORT_1654_COUNT",port_count[1654]);
		     uvm_config_db #(int)::get(null,"","PORT_1655_COUNT",port_count[1655]);
		     uvm_config_db #(int)::get(null,"","PORT_1656_COUNT",port_count[1656]);
		     uvm_config_db #(int)::get(null,"","PORT_1657_COUNT",port_count[1657]);
		     uvm_config_db #(int)::get(null,"","PORT_1658_COUNT",port_count[1658]);
		     uvm_config_db #(int)::get(null,"","PORT_1659_COUNT",port_count[1659]);
		     uvm_config_db #(int)::get(null,"","PORT_1660_COUNT",port_count[1660]);
		     uvm_config_db #(int)::get(null,"","PORT_1661_COUNT",port_count[1661]);
		     uvm_config_db #(int)::get(null,"","PORT_1662_COUNT",port_count[1662]);
		     uvm_config_db #(int)::get(null,"","PORT_1663_COUNT",port_count[1663]);
		     uvm_config_db #(int)::get(null,"","PORT_1664_COUNT",port_count[1664]);
		     uvm_config_db #(int)::get(null,"","PORT_1665_COUNT",port_count[1665]);
		     uvm_config_db #(int)::get(null,"","PORT_1666_COUNT",port_count[1666]);
		     uvm_config_db #(int)::get(null,"","PORT_1667_COUNT",port_count[1667]);
		     uvm_config_db #(int)::get(null,"","PORT_1668_COUNT",port_count[1668]);
		     uvm_config_db #(int)::get(null,"","PORT_1669_COUNT",port_count[1669]);
		     uvm_config_db #(int)::get(null,"","PORT_1670_COUNT",port_count[1670]);
		     uvm_config_db #(int)::get(null,"","PORT_1671_COUNT",port_count[1671]);
		     uvm_config_db #(int)::get(null,"","PORT_1672_COUNT",port_count[1672]);
		     uvm_config_db #(int)::get(null,"","PORT_1673_COUNT",port_count[1673]);
		     uvm_config_db #(int)::get(null,"","PORT_1674_COUNT",port_count[1674]);
		     uvm_config_db #(int)::get(null,"","PORT_1675_COUNT",port_count[1675]);
		     uvm_config_db #(int)::get(null,"","PORT_1676_COUNT",port_count[1676]);
		     uvm_config_db #(int)::get(null,"","PORT_1677_COUNT",port_count[1677]);
		     uvm_config_db #(int)::get(null,"","PORT_1678_COUNT",port_count[1678]);
		     uvm_config_db #(int)::get(null,"","PORT_1679_COUNT",port_count[1679]);
		     uvm_config_db #(int)::get(null,"","PORT_1680_COUNT",port_count[1680]);
		     uvm_config_db #(int)::get(null,"","PORT_1681_COUNT",port_count[1681]);
		     uvm_config_db #(int)::get(null,"","PORT_1682_COUNT",port_count[1682]);
		     uvm_config_db #(int)::get(null,"","PORT_1683_COUNT",port_count[1683]);
		     uvm_config_db #(int)::get(null,"","PORT_1684_COUNT",port_count[1684]);
		     uvm_config_db #(int)::get(null,"","PORT_1685_COUNT",port_count[1685]);
		     uvm_config_db #(int)::get(null,"","PORT_1686_COUNT",port_count[1686]);
		     uvm_config_db #(int)::get(null,"","PORT_1687_COUNT",port_count[1687]);
		     uvm_config_db #(int)::get(null,"","PORT_1688_COUNT",port_count[1688]);
		     uvm_config_db #(int)::get(null,"","PORT_1689_COUNT",port_count[1689]);
		     uvm_config_db #(int)::get(null,"","PORT_1690_COUNT",port_count[1690]);
		     uvm_config_db #(int)::get(null,"","PORT_1691_COUNT",port_count[1691]);
		     uvm_config_db #(int)::get(null,"","PORT_1692_COUNT",port_count[1692]);
		     uvm_config_db #(int)::get(null,"","PORT_1693_COUNT",port_count[1693]);
		     uvm_config_db #(int)::get(null,"","PORT_1694_COUNT",port_count[1694]);
		     uvm_config_db #(int)::get(null,"","PORT_1695_COUNT",port_count[1695]);
		     uvm_config_db #(int)::get(null,"","PORT_1696_COUNT",port_count[1696]);
		     uvm_config_db #(int)::get(null,"","PORT_1697_COUNT",port_count[1697]);
		     uvm_config_db #(int)::get(null,"","PORT_1698_COUNT",port_count[1698]);
		     uvm_config_db #(int)::get(null,"","PORT_1699_COUNT",port_count[1699]);
		     uvm_config_db #(int)::get(null,"","PORT_1700_COUNT",port_count[1700]);
		     uvm_config_db #(int)::get(null,"","PORT_1701_COUNT",port_count[1701]);
		     uvm_config_db #(int)::get(null,"","PORT_1702_COUNT",port_count[1702]);
		     uvm_config_db #(int)::get(null,"","PORT_1703_COUNT",port_count[1703]);
		     uvm_config_db #(int)::get(null,"","PORT_1704_COUNT",port_count[1704]);
		     uvm_config_db #(int)::get(null,"","PORT_1705_COUNT",port_count[1705]);
		     uvm_config_db #(int)::get(null,"","PORT_1706_COUNT",port_count[1706]);
		     uvm_config_db #(int)::get(null,"","PORT_1707_COUNT",port_count[1707]);
		     uvm_config_db #(int)::get(null,"","PORT_1708_COUNT",port_count[1708]);
		     uvm_config_db #(int)::get(null,"","PORT_1709_COUNT",port_count[1709]);
		     uvm_config_db #(int)::get(null,"","PORT_1710_COUNT",port_count[1710]);
		     uvm_config_db #(int)::get(null,"","PORT_1711_COUNT",port_count[1711]);
		     uvm_config_db #(int)::get(null,"","PORT_1712_COUNT",port_count[1712]);
		     uvm_config_db #(int)::get(null,"","PORT_1713_COUNT",port_count[1713]);
		     uvm_config_db #(int)::get(null,"","PORT_1714_COUNT",port_count[1714]);
		     uvm_config_db #(int)::get(null,"","PORT_1715_COUNT",port_count[1715]);
		     uvm_config_db #(int)::get(null,"","PORT_1716_COUNT",port_count[1716]);
		     uvm_config_db #(int)::get(null,"","PORT_1717_COUNT",port_count[1717]);
		     uvm_config_db #(int)::get(null,"","PORT_1718_COUNT",port_count[1718]);
		     uvm_config_db #(int)::get(null,"","PORT_1719_COUNT",port_count[1719]);
		     uvm_config_db #(int)::get(null,"","PORT_1720_COUNT",port_count[1720]);
		     uvm_config_db #(int)::get(null,"","PORT_1721_COUNT",port_count[1721]);
		     uvm_config_db #(int)::get(null,"","PORT_1722_COUNT",port_count[1722]);
		     uvm_config_db #(int)::get(null,"","PORT_1723_COUNT",port_count[1723]);
		     uvm_config_db #(int)::get(null,"","PORT_1724_COUNT",port_count[1724]);
		     uvm_config_db #(int)::get(null,"","PORT_1725_COUNT",port_count[1725]);
		     uvm_config_db #(int)::get(null,"","PORT_1726_COUNT",port_count[1726]);
		     uvm_config_db #(int)::get(null,"","PORT_1727_COUNT",port_count[1727]);
		     uvm_config_db #(int)::get(null,"","PORT_1728_COUNT",port_count[1728]);
		     uvm_config_db #(int)::get(null,"","PORT_1729_COUNT",port_count[1729]);
		     uvm_config_db #(int)::get(null,"","PORT_1730_COUNT",port_count[1730]);
		     uvm_config_db #(int)::get(null,"","PORT_1731_COUNT",port_count[1731]);
		     uvm_config_db #(int)::get(null,"","PORT_1732_COUNT",port_count[1732]);
		     uvm_config_db #(int)::get(null,"","PORT_1733_COUNT",port_count[1733]);
		     uvm_config_db #(int)::get(null,"","PORT_1734_COUNT",port_count[1734]);
		     uvm_config_db #(int)::get(null,"","PORT_1735_COUNT",port_count[1735]);
		     uvm_config_db #(int)::get(null,"","PORT_1736_COUNT",port_count[1736]);
		     uvm_config_db #(int)::get(null,"","PORT_1737_COUNT",port_count[1737]);
		     uvm_config_db #(int)::get(null,"","PORT_1738_COUNT",port_count[1738]);
		     uvm_config_db #(int)::get(null,"","PORT_1739_COUNT",port_count[1739]);
		     uvm_config_db #(int)::get(null,"","PORT_1740_COUNT",port_count[1740]);
		     uvm_config_db #(int)::get(null,"","PORT_1741_COUNT",port_count[1741]);
		     uvm_config_db #(int)::get(null,"","PORT_1742_COUNT",port_count[1742]);
		     uvm_config_db #(int)::get(null,"","PORT_1743_COUNT",port_count[1743]);
		     uvm_config_db #(int)::get(null,"","PORT_1744_COUNT",port_count[1744]);
		     uvm_config_db #(int)::get(null,"","PORT_1745_COUNT",port_count[1745]);
		     uvm_config_db #(int)::get(null,"","PORT_1746_COUNT",port_count[1746]);
		     uvm_config_db #(int)::get(null,"","PORT_1747_COUNT",port_count[1747]);
		     uvm_config_db #(int)::get(null,"","PORT_1748_COUNT",port_count[1748]);
		     uvm_config_db #(int)::get(null,"","PORT_1749_COUNT",port_count[1749]);
		     uvm_config_db #(int)::get(null,"","PORT_1750_COUNT",port_count[1750]);
		     uvm_config_db #(int)::get(null,"","PORT_1751_COUNT",port_count[1751]);
		     uvm_config_db #(int)::get(null,"","PORT_1752_COUNT",port_count[1752]);
		     uvm_config_db #(int)::get(null,"","PORT_1753_COUNT",port_count[1753]);
		     uvm_config_db #(int)::get(null,"","PORT_1754_COUNT",port_count[1754]);
		     uvm_config_db #(int)::get(null,"","PORT_1755_COUNT",port_count[1755]);
		     uvm_config_db #(int)::get(null,"","PORT_1756_COUNT",port_count[1756]);
		     uvm_config_db #(int)::get(null,"","PORT_1757_COUNT",port_count[1757]);
		     uvm_config_db #(int)::get(null,"","PORT_1758_COUNT",port_count[1758]);
		     uvm_config_db #(int)::get(null,"","PORT_1759_COUNT",port_count[1759]);
		     uvm_config_db #(int)::get(null,"","PORT_1760_COUNT",port_count[1760]);
		     uvm_config_db #(int)::get(null,"","PORT_1761_COUNT",port_count[1761]);
		     uvm_config_db #(int)::get(null,"","PORT_1762_COUNT",port_count[1762]);
		     uvm_config_db #(int)::get(null,"","PORT_1763_COUNT",port_count[1763]);
		     uvm_config_db #(int)::get(null,"","PORT_1764_COUNT",port_count[1764]);
		     uvm_config_db #(int)::get(null,"","PORT_1765_COUNT",port_count[1765]);
		     uvm_config_db #(int)::get(null,"","PORT_1766_COUNT",port_count[1766]);
		     uvm_config_db #(int)::get(null,"","PORT_1767_COUNT",port_count[1767]);
		     uvm_config_db #(int)::get(null,"","PORT_1768_COUNT",port_count[1768]);
		     uvm_config_db #(int)::get(null,"","PORT_1769_COUNT",port_count[1769]);
		     uvm_config_db #(int)::get(null,"","PORT_1770_COUNT",port_count[1770]);
		     uvm_config_db #(int)::get(null,"","PORT_1771_COUNT",port_count[1771]);
		     uvm_config_db #(int)::get(null,"","PORT_1772_COUNT",port_count[1772]);
		     uvm_config_db #(int)::get(null,"","PORT_1773_COUNT",port_count[1773]);
		     uvm_config_db #(int)::get(null,"","PORT_1774_COUNT",port_count[1774]);
		     uvm_config_db #(int)::get(null,"","PORT_1775_COUNT",port_count[1775]);
		     uvm_config_db #(int)::get(null,"","PORT_1776_COUNT",port_count[1776]);
		     uvm_config_db #(int)::get(null,"","PORT_1777_COUNT",port_count[1777]);
		     uvm_config_db #(int)::get(null,"","PORT_1778_COUNT",port_count[1778]);
		     uvm_config_db #(int)::get(null,"","PORT_1779_COUNT",port_count[1779]);
		     uvm_config_db #(int)::get(null,"","PORT_1780_COUNT",port_count[1780]);
		     uvm_config_db #(int)::get(null,"","PORT_1781_COUNT",port_count[1781]);
		     uvm_config_db #(int)::get(null,"","PORT_1782_COUNT",port_count[1782]);
		     uvm_config_db #(int)::get(null,"","PORT_1783_COUNT",port_count[1783]);
		     uvm_config_db #(int)::get(null,"","PORT_1784_COUNT",port_count[1784]);
		     uvm_config_db #(int)::get(null,"","PORT_1785_COUNT",port_count[1785]);
		     uvm_config_db #(int)::get(null,"","PORT_1786_COUNT",port_count[1786]);
		     uvm_config_db #(int)::get(null,"","PORT_1787_COUNT",port_count[1787]);
		     uvm_config_db #(int)::get(null,"","PORT_1788_COUNT",port_count[1788]);
		     uvm_config_db #(int)::get(null,"","PORT_1789_COUNT",port_count[1789]);
		     uvm_config_db #(int)::get(null,"","PORT_1790_COUNT",port_count[1790]);
		     uvm_config_db #(int)::get(null,"","PORT_1791_COUNT",port_count[1791]);
		     uvm_config_db #(int)::get(null,"","PORT_1792_COUNT",port_count[1792]);
		     uvm_config_db #(int)::get(null,"","PORT_1793_COUNT",port_count[1793]);
		     uvm_config_db #(int)::get(null,"","PORT_1794_COUNT",port_count[1794]);
		     uvm_config_db #(int)::get(null,"","PORT_1795_COUNT",port_count[1795]);
		     uvm_config_db #(int)::get(null,"","PORT_1796_COUNT",port_count[1796]);
		     uvm_config_db #(int)::get(null,"","PORT_1797_COUNT",port_count[1797]);
		     uvm_config_db #(int)::get(null,"","PORT_1798_COUNT",port_count[1798]);
		     uvm_config_db #(int)::get(null,"","PORT_1799_COUNT",port_count[1799]);
		     uvm_config_db #(int)::get(null,"","PORT_1800_COUNT",port_count[1800]);
		     uvm_config_db #(int)::get(null,"","PORT_1801_COUNT",port_count[1801]);
		     uvm_config_db #(int)::get(null,"","PORT_1802_COUNT",port_count[1802]);
		     uvm_config_db #(int)::get(null,"","PORT_1803_COUNT",port_count[1803]);
		     uvm_config_db #(int)::get(null,"","PORT_1804_COUNT",port_count[1804]);
		     uvm_config_db #(int)::get(null,"","PORT_1805_COUNT",port_count[1805]);
		     uvm_config_db #(int)::get(null,"","PORT_1806_COUNT",port_count[1806]);
		     uvm_config_db #(int)::get(null,"","PORT_1807_COUNT",port_count[1807]);
		     uvm_config_db #(int)::get(null,"","PORT_1808_COUNT",port_count[1808]);
		     uvm_config_db #(int)::get(null,"","PORT_1809_COUNT",port_count[1809]);
		     uvm_config_db #(int)::get(null,"","PORT_1810_COUNT",port_count[1810]);
		     uvm_config_db #(int)::get(null,"","PORT_1811_COUNT",port_count[1811]);
		     uvm_config_db #(int)::get(null,"","PORT_1812_COUNT",port_count[1812]);
		     uvm_config_db #(int)::get(null,"","PORT_1813_COUNT",port_count[1813]);
		     uvm_config_db #(int)::get(null,"","PORT_1814_COUNT",port_count[1814]);
		     uvm_config_db #(int)::get(null,"","PORT_1815_COUNT",port_count[1815]);
		     uvm_config_db #(int)::get(null,"","PORT_1816_COUNT",port_count[1816]);
		     uvm_config_db #(int)::get(null,"","PORT_1817_COUNT",port_count[1817]);
		     uvm_config_db #(int)::get(null,"","PORT_1818_COUNT",port_count[1818]);
		     uvm_config_db #(int)::get(null,"","PORT_1819_COUNT",port_count[1819]);
		     uvm_config_db #(int)::get(null,"","PORT_1820_COUNT",port_count[1820]);
		     uvm_config_db #(int)::get(null,"","PORT_1821_COUNT",port_count[1821]);
		     uvm_config_db #(int)::get(null,"","PORT_1822_COUNT",port_count[1822]);
		     uvm_config_db #(int)::get(null,"","PORT_1823_COUNT",port_count[1823]);
		     uvm_config_db #(int)::get(null,"","PORT_1824_COUNT",port_count[1824]);
		     uvm_config_db #(int)::get(null,"","PORT_1825_COUNT",port_count[1825]);
		     uvm_config_db #(int)::get(null,"","PORT_1826_COUNT",port_count[1826]);
		     uvm_config_db #(int)::get(null,"","PORT_1827_COUNT",port_count[1827]);
		     uvm_config_db #(int)::get(null,"","PORT_1828_COUNT",port_count[1828]);
		     uvm_config_db #(int)::get(null,"","PORT_1829_COUNT",port_count[1829]);
		     uvm_config_db #(int)::get(null,"","PORT_1830_COUNT",port_count[1830]);
		     uvm_config_db #(int)::get(null,"","PORT_1831_COUNT",port_count[1831]);
		     uvm_config_db #(int)::get(null,"","PORT_1832_COUNT",port_count[1832]);
		     uvm_config_db #(int)::get(null,"","PORT_1833_COUNT",port_count[1833]);
		     uvm_config_db #(int)::get(null,"","PORT_1834_COUNT",port_count[1834]);
		     uvm_config_db #(int)::get(null,"","PORT_1835_COUNT",port_count[1835]);
		     uvm_config_db #(int)::get(null,"","PORT_1836_COUNT",port_count[1836]);
		     uvm_config_db #(int)::get(null,"","PORT_1837_COUNT",port_count[1837]);
		     uvm_config_db #(int)::get(null,"","PORT_1838_COUNT",port_count[1838]);
		     uvm_config_db #(int)::get(null,"","PORT_1839_COUNT",port_count[1839]);
		     uvm_config_db #(int)::get(null,"","PORT_1840_COUNT",port_count[1840]);
		     uvm_config_db #(int)::get(null,"","PORT_1841_COUNT",port_count[1841]);
		     uvm_config_db #(int)::get(null,"","PORT_1842_COUNT",port_count[1842]);
		     uvm_config_db #(int)::get(null,"","PORT_1843_COUNT",port_count[1843]);
		     uvm_config_db #(int)::get(null,"","PORT_1844_COUNT",port_count[1844]);
		     uvm_config_db #(int)::get(null,"","PORT_1845_COUNT",port_count[1845]);
		     uvm_config_db #(int)::get(null,"","PORT_1846_COUNT",port_count[1846]);
		     uvm_config_db #(int)::get(null,"","PORT_1847_COUNT",port_count[1847]);
		     uvm_config_db #(int)::get(null,"","PORT_1848_COUNT",port_count[1848]);
		     uvm_config_db #(int)::get(null,"","PORT_1849_COUNT",port_count[1849]);
		     uvm_config_db #(int)::get(null,"","PORT_1850_COUNT",port_count[1850]);
		     uvm_config_db #(int)::get(null,"","PORT_1851_COUNT",port_count[1851]);
		     uvm_config_db #(int)::get(null,"","PORT_1852_COUNT",port_count[1852]);
		     uvm_config_db #(int)::get(null,"","PORT_1853_COUNT",port_count[1853]);
		     uvm_config_db #(int)::get(null,"","PORT_1854_COUNT",port_count[1854]);
		     uvm_config_db #(int)::get(null,"","PORT_1855_COUNT",port_count[1855]);
		     uvm_config_db #(int)::get(null,"","PORT_1856_COUNT",port_count[1856]);
		     uvm_config_db #(int)::get(null,"","PORT_1857_COUNT",port_count[1857]);
		     uvm_config_db #(int)::get(null,"","PORT_1858_COUNT",port_count[1858]);
		     uvm_config_db #(int)::get(null,"","PORT_1859_COUNT",port_count[1859]);
		     uvm_config_db #(int)::get(null,"","PORT_1860_COUNT",port_count[1860]);
		     uvm_config_db #(int)::get(null,"","PORT_1861_COUNT",port_count[1861]);
		     uvm_config_db #(int)::get(null,"","PORT_1862_COUNT",port_count[1862]);
		     uvm_config_db #(int)::get(null,"","PORT_1863_COUNT",port_count[1863]);
		     uvm_config_db #(int)::get(null,"","PORT_1864_COUNT",port_count[1864]);
		     uvm_config_db #(int)::get(null,"","PORT_1865_COUNT",port_count[1865]);
		     uvm_config_db #(int)::get(null,"","PORT_1866_COUNT",port_count[1866]);
		     uvm_config_db #(int)::get(null,"","PORT_1867_COUNT",port_count[1867]);
		     uvm_config_db #(int)::get(null,"","PORT_1868_COUNT",port_count[1868]);
		     uvm_config_db #(int)::get(null,"","PORT_1869_COUNT",port_count[1869]);
		     uvm_config_db #(int)::get(null,"","PORT_1870_COUNT",port_count[1870]);
		     uvm_config_db #(int)::get(null,"","PORT_1871_COUNT",port_count[1871]);
		     uvm_config_db #(int)::get(null,"","PORT_1872_COUNT",port_count[1872]);
		     uvm_config_db #(int)::get(null,"","PORT_1873_COUNT",port_count[1873]);
		     uvm_config_db #(int)::get(null,"","PORT_1874_COUNT",port_count[1874]);
		     uvm_config_db #(int)::get(null,"","PORT_1875_COUNT",port_count[1875]);
		     uvm_config_db #(int)::get(null,"","PORT_1876_COUNT",port_count[1876]);
		     uvm_config_db #(int)::get(null,"","PORT_1877_COUNT",port_count[1877]);
		     uvm_config_db #(int)::get(null,"","PORT_1878_COUNT",port_count[1878]);
		     uvm_config_db #(int)::get(null,"","PORT_1879_COUNT",port_count[1879]);
		     uvm_config_db #(int)::get(null,"","PORT_1880_COUNT",port_count[1880]);
		     uvm_config_db #(int)::get(null,"","PORT_1881_COUNT",port_count[1881]);
		     uvm_config_db #(int)::get(null,"","PORT_1882_COUNT",port_count[1882]);
		     uvm_config_db #(int)::get(null,"","PORT_1883_COUNT",port_count[1883]);
		     uvm_config_db #(int)::get(null,"","PORT_1884_COUNT",port_count[1884]);
		     uvm_config_db #(int)::get(null,"","PORT_1885_COUNT",port_count[1885]);
		     uvm_config_db #(int)::get(null,"","PORT_1886_COUNT",port_count[1886]);
		     uvm_config_db #(int)::get(null,"","PORT_1887_COUNT",port_count[1887]);
		     uvm_config_db #(int)::get(null,"","PORT_1888_COUNT",port_count[1888]);
		     uvm_config_db #(int)::get(null,"","PORT_1889_COUNT",port_count[1889]);
		     uvm_config_db #(int)::get(null,"","PORT_1890_COUNT",port_count[1890]);
		     uvm_config_db #(int)::get(null,"","PORT_1891_COUNT",port_count[1891]);
		     uvm_config_db #(int)::get(null,"","PORT_1892_COUNT",port_count[1892]);
		     uvm_config_db #(int)::get(null,"","PORT_1893_COUNT",port_count[1893]);
		     uvm_config_db #(int)::get(null,"","PORT_1894_COUNT",port_count[1894]);
		     uvm_config_db #(int)::get(null,"","PORT_1895_COUNT",port_count[1895]);
		     uvm_config_db #(int)::get(null,"","PORT_1896_COUNT",port_count[1896]);
		     uvm_config_db #(int)::get(null,"","PORT_1897_COUNT",port_count[1897]);
		     uvm_config_db #(int)::get(null,"","PORT_1898_COUNT",port_count[1898]);
		     uvm_config_db #(int)::get(null,"","PORT_1899_COUNT",port_count[1899]);
		     uvm_config_db #(int)::get(null,"","PORT_1900_COUNT",port_count[1900]);
		     uvm_config_db #(int)::get(null,"","PORT_1901_COUNT",port_count[1901]);
		     uvm_config_db #(int)::get(null,"","PORT_1902_COUNT",port_count[1902]);
		     uvm_config_db #(int)::get(null,"","PORT_1903_COUNT",port_count[1903]);
		     uvm_config_db #(int)::get(null,"","PORT_1904_COUNT",port_count[1904]);
		     uvm_config_db #(int)::get(null,"","PORT_1905_COUNT",port_count[1905]);
		     uvm_config_db #(int)::get(null,"","PORT_1906_COUNT",port_count[1906]);
		     uvm_config_db #(int)::get(null,"","PORT_1907_COUNT",port_count[1907]);
		     uvm_config_db #(int)::get(null,"","PORT_1908_COUNT",port_count[1908]);
		     uvm_config_db #(int)::get(null,"","PORT_1909_COUNT",port_count[1909]);
		     uvm_config_db #(int)::get(null,"","PORT_1910_COUNT",port_count[1910]);
		     uvm_config_db #(int)::get(null,"","PORT_1911_COUNT",port_count[1911]);
		     uvm_config_db #(int)::get(null,"","PORT_1912_COUNT",port_count[1912]);
		     uvm_config_db #(int)::get(null,"","PORT_1913_COUNT",port_count[1913]);
		     uvm_config_db #(int)::get(null,"","PORT_1914_COUNT",port_count[1914]);
		     uvm_config_db #(int)::get(null,"","PORT_1915_COUNT",port_count[1915]);
		     uvm_config_db #(int)::get(null,"","PORT_1916_COUNT",port_count[1916]);
		     uvm_config_db #(int)::get(null,"","PORT_1917_COUNT",port_count[1917]);
		     uvm_config_db #(int)::get(null,"","PORT_1918_COUNT",port_count[1918]);
		     uvm_config_db #(int)::get(null,"","PORT_1919_COUNT",port_count[1919]);
		     uvm_config_db #(int)::get(null,"","PORT_1920_COUNT",port_count[1920]);
		     uvm_config_db #(int)::get(null,"","PORT_1921_COUNT",port_count[1921]);
		     uvm_config_db #(int)::get(null,"","PORT_1922_COUNT",port_count[1922]);
		     uvm_config_db #(int)::get(null,"","PORT_1923_COUNT",port_count[1923]);
		     uvm_config_db #(int)::get(null,"","PORT_1924_COUNT",port_count[1924]);
		     uvm_config_db #(int)::get(null,"","PORT_1925_COUNT",port_count[1925]);
		     uvm_config_db #(int)::get(null,"","PORT_1926_COUNT",port_count[1926]);
		     uvm_config_db #(int)::get(null,"","PORT_1927_COUNT",port_count[1927]);
		     uvm_config_db #(int)::get(null,"","PORT_1928_COUNT",port_count[1928]);
		     uvm_config_db #(int)::get(null,"","PORT_1929_COUNT",port_count[1929]);
		     uvm_config_db #(int)::get(null,"","PORT_1930_COUNT",port_count[1930]);
		     uvm_config_db #(int)::get(null,"","PORT_1931_COUNT",port_count[1931]);
		     uvm_config_db #(int)::get(null,"","PORT_1932_COUNT",port_count[1932]);
		     uvm_config_db #(int)::get(null,"","PORT_1933_COUNT",port_count[1933]);
		     uvm_config_db #(int)::get(null,"","PORT_1934_COUNT",port_count[1934]);
		     uvm_config_db #(int)::get(null,"","PORT_1935_COUNT",port_count[1935]);
		     uvm_config_db #(int)::get(null,"","PORT_1936_COUNT",port_count[1936]);
		     uvm_config_db #(int)::get(null,"","PORT_1937_COUNT",port_count[1937]);
		     uvm_config_db #(int)::get(null,"","PORT_1938_COUNT",port_count[1938]);
		     uvm_config_db #(int)::get(null,"","PORT_1939_COUNT",port_count[1939]);
		     uvm_config_db #(int)::get(null,"","PORT_1940_COUNT",port_count[1940]);
		     uvm_config_db #(int)::get(null,"","PORT_1941_COUNT",port_count[1941]);
		     uvm_config_db #(int)::get(null,"","PORT_1942_COUNT",port_count[1942]);
		     uvm_config_db #(int)::get(null,"","PORT_1943_COUNT",port_count[1943]);
		     uvm_config_db #(int)::get(null,"","PORT_1944_COUNT",port_count[1944]);
		     uvm_config_db #(int)::get(null,"","PORT_1945_COUNT",port_count[1945]);
		     uvm_config_db #(int)::get(null,"","PORT_1946_COUNT",port_count[1946]);
		     uvm_config_db #(int)::get(null,"","PORT_1947_COUNT",port_count[1947]);
		     uvm_config_db #(int)::get(null,"","PORT_1948_COUNT",port_count[1948]);
		     uvm_config_db #(int)::get(null,"","PORT_1949_COUNT",port_count[1949]);
		     uvm_config_db #(int)::get(null,"","PORT_1950_COUNT",port_count[1950]);
		     uvm_config_db #(int)::get(null,"","PORT_1951_COUNT",port_count[1951]);
		     uvm_config_db #(int)::get(null,"","PORT_1952_COUNT",port_count[1952]);
		     uvm_config_db #(int)::get(null,"","PORT_1953_COUNT",port_count[1953]);
		     uvm_config_db #(int)::get(null,"","PORT_1954_COUNT",port_count[1954]);
		     uvm_config_db #(int)::get(null,"","PORT_1955_COUNT",port_count[1955]);
		     uvm_config_db #(int)::get(null,"","PORT_1956_COUNT",port_count[1956]);
		     uvm_config_db #(int)::get(null,"","PORT_1957_COUNT",port_count[1957]);
		     uvm_config_db #(int)::get(null,"","PORT_1958_COUNT",port_count[1958]);
		     uvm_config_db #(int)::get(null,"","PORT_1959_COUNT",port_count[1959]);
		     uvm_config_db #(int)::get(null,"","PORT_1960_COUNT",port_count[1960]);
		     uvm_config_db #(int)::get(null,"","PORT_1961_COUNT",port_count[1961]);
		     uvm_config_db #(int)::get(null,"","PORT_1962_COUNT",port_count[1962]);
		     uvm_config_db #(int)::get(null,"","PORT_1963_COUNT",port_count[1963]);
		     uvm_config_db #(int)::get(null,"","PORT_1964_COUNT",port_count[1964]);
		     uvm_config_db #(int)::get(null,"","PORT_1965_COUNT",port_count[1965]);
		     uvm_config_db #(int)::get(null,"","PORT_1966_COUNT",port_count[1966]);
		     uvm_config_db #(int)::get(null,"","PORT_1967_COUNT",port_count[1967]);
		     uvm_config_db #(int)::get(null,"","PORT_1968_COUNT",port_count[1968]);
		     uvm_config_db #(int)::get(null,"","PORT_1969_COUNT",port_count[1969]);
		     uvm_config_db #(int)::get(null,"","PORT_1970_COUNT",port_count[1970]);
		     uvm_config_db #(int)::get(null,"","PORT_1971_COUNT",port_count[1971]);
		     uvm_config_db #(int)::get(null,"","PORT_1972_COUNT",port_count[1972]);
		     uvm_config_db #(int)::get(null,"","PORT_1973_COUNT",port_count[1973]);
		     uvm_config_db #(int)::get(null,"","PORT_1974_COUNT",port_count[1974]);
		     uvm_config_db #(int)::get(null,"","PORT_1975_COUNT",port_count[1975]);
		     uvm_config_db #(int)::get(null,"","PORT_1976_COUNT",port_count[1976]);
		     uvm_config_db #(int)::get(null,"","PORT_1977_COUNT",port_count[1977]);
		     uvm_config_db #(int)::get(null,"","PORT_1978_COUNT",port_count[1978]);
		     uvm_config_db #(int)::get(null,"","PORT_1979_COUNT",port_count[1979]);
		     uvm_config_db #(int)::get(null,"","PORT_1980_COUNT",port_count[1980]);
		     uvm_config_db #(int)::get(null,"","PORT_1981_COUNT",port_count[1981]);
		     uvm_config_db #(int)::get(null,"","PORT_1982_COUNT",port_count[1982]);
		     uvm_config_db #(int)::get(null,"","PORT_1983_COUNT",port_count[1983]);
		     uvm_config_db #(int)::get(null,"","PORT_1984_COUNT",port_count[1984]);
		     uvm_config_db #(int)::get(null,"","PORT_1985_COUNT",port_count[1985]);
		     uvm_config_db #(int)::get(null,"","PORT_1986_COUNT",port_count[1986]);
		     uvm_config_db #(int)::get(null,"","PORT_1987_COUNT",port_count[1987]);
		     uvm_config_db #(int)::get(null,"","PORT_1988_COUNT",port_count[1988]);
		     uvm_config_db #(int)::get(null,"","PORT_1989_COUNT",port_count[1989]);
		     uvm_config_db #(int)::get(null,"","PORT_1990_COUNT",port_count[1990]);
		     uvm_config_db #(int)::get(null,"","PORT_1991_COUNT",port_count[1991]);
		     uvm_config_db #(int)::get(null,"","PORT_1992_COUNT",port_count[1992]);
		     uvm_config_db #(int)::get(null,"","PORT_1993_COUNT",port_count[1993]);
		     uvm_config_db #(int)::get(null,"","PORT_1994_COUNT",port_count[1994]);
		     uvm_config_db #(int)::get(null,"","PORT_1995_COUNT",port_count[1995]);
		     uvm_config_db #(int)::get(null,"","PORT_1996_COUNT",port_count[1996]);
		     uvm_config_db #(int)::get(null,"","PORT_1997_COUNT",port_count[1997]);
		     uvm_config_db #(int)::get(null,"","PORT_1998_COUNT",port_count[1998]);
		     uvm_config_db #(int)::get(null,"","PORT_1999_COUNT",port_count[1999]);
		     uvm_config_db #(int)::get(null,"","PORT_2000_COUNT",port_count[2000]);
		     uvm_config_db #(int)::get(null,"","PORT_2001_COUNT",port_count[2001]);
		     uvm_config_db #(int)::get(null,"","PORT_2002_COUNT",port_count[2002]);
		     uvm_config_db #(int)::get(null,"","PORT_2003_COUNT",port_count[2003]);
		     uvm_config_db #(int)::get(null,"","PORT_2004_COUNT",port_count[2004]);
		     uvm_config_db #(int)::get(null,"","PORT_2005_COUNT",port_count[2005]);
		     uvm_config_db #(int)::get(null,"","PORT_2006_COUNT",port_count[2006]);
		     uvm_config_db #(int)::get(null,"","PORT_2007_COUNT",port_count[2007]);
		     uvm_config_db #(int)::get(null,"","PORT_2008_COUNT",port_count[2008]);
		     uvm_config_db #(int)::get(null,"","PORT_2009_COUNT",port_count[2009]);
		     uvm_config_db #(int)::get(null,"","PORT_2010_COUNT",port_count[2010]);
		     uvm_config_db #(int)::get(null,"","PORT_2011_COUNT",port_count[2011]);
		     uvm_config_db #(int)::get(null,"","PORT_2012_COUNT",port_count[2012]);
		     uvm_config_db #(int)::get(null,"","PORT_2013_COUNT",port_count[2013]);
		     uvm_config_db #(int)::get(null,"","PORT_2014_COUNT",port_count[2014]);
		     uvm_config_db #(int)::get(null,"","PORT_2015_COUNT",port_count[2015]);
		     uvm_config_db #(int)::get(null,"","PORT_2016_COUNT",port_count[2016]);
		     uvm_config_db #(int)::get(null,"","PORT_2017_COUNT",port_count[2017]);
		     uvm_config_db #(int)::get(null,"","PORT_2018_COUNT",port_count[2018]);
		     uvm_config_db #(int)::get(null,"","PORT_2019_COUNT",port_count[2019]);
		     uvm_config_db #(int)::get(null,"","PORT_2020_COUNT",port_count[2020]);
		     uvm_config_db #(int)::get(null,"","PORT_2021_COUNT",port_count[2021]);
		     uvm_config_db #(int)::get(null,"","PORT_2022_COUNT",port_count[2022]);
		     uvm_config_db #(int)::get(null,"","PORT_2023_COUNT",port_count[2023]);
		     uvm_config_db #(int)::get(null,"","PORT_2024_COUNT",port_count[2024]);
		     uvm_config_db #(int)::get(null,"","PORT_2025_COUNT",port_count[2025]);
		     uvm_config_db #(int)::get(null,"","PORT_2026_COUNT",port_count[2026]);
		     uvm_config_db #(int)::get(null,"","PORT_2027_COUNT",port_count[2027]);
		     uvm_config_db #(int)::get(null,"","PORT_2028_COUNT",port_count[2028]);
		     uvm_config_db #(int)::get(null,"","PORT_2029_COUNT",port_count[2029]);
		     uvm_config_db #(int)::get(null,"","PORT_2030_COUNT",port_count[2030]);
		     uvm_config_db #(int)::get(null,"","PORT_2031_COUNT",port_count[2031]);
		     uvm_config_db #(int)::get(null,"","PORT_2032_COUNT",port_count[2032]);
		     uvm_config_db #(int)::get(null,"","PORT_2033_COUNT",port_count[2033]);
		     uvm_config_db #(int)::get(null,"","PORT_2034_COUNT",port_count[2034]);
		     uvm_config_db #(int)::get(null,"","PORT_2035_COUNT",port_count[2035]);
		     uvm_config_db #(int)::get(null,"","PORT_2036_COUNT",port_count[2036]);
		     uvm_config_db #(int)::get(null,"","PORT_2037_COUNT",port_count[2037]);
		     uvm_config_db #(int)::get(null,"","PORT_2038_COUNT",port_count[2038]);
		     uvm_config_db #(int)::get(null,"","PORT_2039_COUNT",port_count[2039]);
		     uvm_config_db #(int)::get(null,"","PORT_2040_COUNT",port_count[2040]);
		     uvm_config_db #(int)::get(null,"","PORT_2041_COUNT",port_count[2041]);
		     uvm_config_db #(int)::get(null,"","PORT_2042_COUNT",port_count[2042]);
		     uvm_config_db #(int)::get(null,"","PORT_2043_COUNT",port_count[2043]);
		     uvm_config_db #(int)::get(null,"","PORT_2044_COUNT",port_count[2044]);
		     uvm_config_db #(int)::get(null,"","PORT_2045_COUNT",port_count[2045]);
		     uvm_config_db #(int)::get(null,"","PORT_2046_COUNT",port_count[2046]);
		     uvm_config_db #(int)::get(null,"","PORT_2047_COUNT",port_count[2047]);
         `endif
      packet_count_check(port_count[0],env.pf_vf_mux_scbd_0.packet_count,0);
      packet_count_check(port_count[1],env.pf_vf_mux_scbd_1.packet_count,1);
      packet_count_check(port_count[2],env.pf_vf_mux_scbd_2.packet_count,2);
      packet_count_check(port_count[3],env.pf_vf_mux_scbd_3.packet_count,3);
      packet_count_check(port_count[4],env.pf_vf_mux_scbd_4.packet_count,4);
      packet_count_check(port_count[5],env.pf_vf_mux_scbd_5.packet_count,5);
      packet_count_check(port_count[6],env.pf_vf_mux_scbd_6.packet_count,6);
      packet_count_check(port_count[7],env.pf_vf_mux_scbd_7.packet_count,7);
      packet_count_check(port_count[8],env.pf_vf_mux_scbd_8.packet_count,8);
      packet_count_check(port_count[9],env.pf_vf_mux_scbd_9.packet_count,9);
      packet_count_check(port_count[10],env.pf_vf_mux_scbd_10.packet_count,10);
      packet_count_check(port_count[11],env.pf_vf_mux_scbd_11.packet_count,11);
      packet_count_check(port_count[12],env.pf_vf_mux_scbd_12.packet_count,12);
      packet_count_check(port_count[13],env.pf_vf_mux_scbd_13.packet_count,13);
      packet_count_check(port_count[14],env.pf_vf_mux_scbd_14.packet_count,14);
      packet_count_check(port_count[15],env.pf_vf_mux_scbd_15.packet_count,15);
      `ifdef TB_CONFIG_2
      packet_count_check(port_count[16],env.pf_vf_mux_scbd_16.packet_count,16);
      packet_count_check(port_count[17],env.pf_vf_mux_scbd_17.packet_count,17);
      packet_count_check(port_count[18],env.pf_vf_mux_scbd_18.packet_count,18);
      packet_count_check(port_count[19],env.pf_vf_mux_scbd_19.packet_count,19);
      packet_count_check(port_count[20],env.pf_vf_mux_scbd_20.packet_count,20);
      packet_count_check(port_count[21],env.pf_vf_mux_scbd_21.packet_count,21);
      packet_count_check(port_count[22],env.pf_vf_mux_scbd_22.packet_count,22);
      packet_count_check(port_count[23],env.pf_vf_mux_scbd_23.packet_count,23);
      `elsif TB_CONFIG_3
      packet_count_check(port_count[16],env.pf_vf_mux_scbd_16.packet_count,16);
      packet_count_check(port_count[17],env.pf_vf_mux_scbd_17.packet_count,17);
      packet_count_check(port_count[18],env.pf_vf_mux_scbd_18.packet_count,18);
      packet_count_check(port_count[19],env.pf_vf_mux_scbd_19.packet_count,19);
      packet_count_check(port_count[20],env.pf_vf_mux_scbd_20.packet_count,20);
      packet_count_check(port_count[21],env.pf_vf_mux_scbd_21.packet_count,21);
      packet_count_check(port_count[22],env.pf_vf_mux_scbd_22.packet_count,22);
      packet_count_check(port_count[23],env.pf_vf_mux_scbd_23.packet_count,23);
      packet_count_check(port_count[24],env.pf_vf_mux_scbd_24.packet_count,24);
      packet_count_check(port_count[25],env.pf_vf_mux_scbd_25.packet_count,25);
      packet_count_check(port_count[26],env.pf_vf_mux_scbd_26.packet_count,26);
      packet_count_check(port_count[27],env.pf_vf_mux_scbd_27.packet_count,27);
      packet_count_check(port_count[28],env.pf_vf_mux_scbd_28.packet_count,28);
      packet_count_check(port_count[29],env.pf_vf_mux_scbd_29.packet_count,29);
      packet_count_check(port_count[30],env.pf_vf_mux_scbd_30.packet_count,30);
      packet_count_check(port_count[31],env.pf_vf_mux_scbd_31.packet_count,31);
      `elsif TB_CONFIG_4
      packet_count_check(port_count[16],env.pf_vf_mux_scbd_16.packet_count,16);
      packet_count_check(port_count[17],env.pf_vf_mux_scbd_17.packet_count,17);
      packet_count_check(port_count[18],env.pf_vf_mux_scbd_18.packet_count,18);
      packet_count_check(port_count[19],env.pf_vf_mux_scbd_19.packet_count,19);
      packet_count_check(port_count[20],env.pf_vf_mux_scbd_20.packet_count,20);
      packet_count_check(port_count[21],env.pf_vf_mux_scbd_21.packet_count,21);
      packet_count_check(port_count[22],env.pf_vf_mux_scbd_22.packet_count,22);
      packet_count_check(port_count[23],env.pf_vf_mux_scbd_23.packet_count,23);
      packet_count_check(port_count[24],env.pf_vf_mux_scbd_24.packet_count,24);
      packet_count_check(port_count[25],env.pf_vf_mux_scbd_25.packet_count,25);
      packet_count_check(port_count[26],env.pf_vf_mux_scbd_26.packet_count,26);
      packet_count_check(port_count[27],env.pf_vf_mux_scbd_27.packet_count,27);
      packet_count_check(port_count[28],env.pf_vf_mux_scbd_28.packet_count,28);
      packet_count_check(port_count[29],env.pf_vf_mux_scbd_29.packet_count,29);
      packet_count_check(port_count[30],env.pf_vf_mux_scbd_30.packet_count,30);
      packet_count_check(port_count[31],env.pf_vf_mux_scbd_31.packet_count,31);
      packet_count_check(port_count[32],env.pf_vf_mux_scbd_32.packet_count,32);
      packet_count_check(port_count[33],env.pf_vf_mux_scbd_33.packet_count,33);
      packet_count_check(port_count[34],env.pf_vf_mux_scbd_34.packet_count,34);
      packet_count_check(port_count[35],env.pf_vf_mux_scbd_35.packet_count,35);
      packet_count_check(port_count[36],env.pf_vf_mux_scbd_36.packet_count,36);
      packet_count_check(port_count[37],env.pf_vf_mux_scbd_37.packet_count,37);
      packet_count_check(port_count[38],env.pf_vf_mux_scbd_38.packet_count,38);
      packet_count_check(port_count[39],env.pf_vf_mux_scbd_39.packet_count,39);
      packet_count_check(port_count[40],env.pf_vf_mux_scbd_40.packet_count,40);
      packet_count_check(port_count[41],env.pf_vf_mux_scbd_41.packet_count,41);
      packet_count_check(port_count[42],env.pf_vf_mux_scbd_42.packet_count,42);
      packet_count_check(port_count[43],env.pf_vf_mux_scbd_43.packet_count,43);
      packet_count_check(port_count[44],env.pf_vf_mux_scbd_44.packet_count,44);
      packet_count_check(port_count[45],env.pf_vf_mux_scbd_45.packet_count,45);
      packet_count_check(port_count[46],env.pf_vf_mux_scbd_46.packet_count,46);
      packet_count_check(port_count[47],env.pf_vf_mux_scbd_47.packet_count,47);
      packet_count_check(port_count[48],env.pf_vf_mux_scbd_48.packet_count,48);
      packet_count_check(port_count[49],env.pf_vf_mux_scbd_49.packet_count,49);
      packet_count_check(port_count[50],env.pf_vf_mux_scbd_50.packet_count,50);
      packet_count_check(port_count[51],env.pf_vf_mux_scbd_51.packet_count,51);
      packet_count_check(port_count[52],env.pf_vf_mux_scbd_52.packet_count,52);
      packet_count_check(port_count[53],env.pf_vf_mux_scbd_53.packet_count,53);
      packet_count_check(port_count[54],env.pf_vf_mux_scbd_54.packet_count,54);
      packet_count_check(port_count[55],env.pf_vf_mux_scbd_55.packet_count,55);
      packet_count_check(port_count[56],env.pf_vf_mux_scbd_56.packet_count,56);
      packet_count_check(port_count[57],env.pf_vf_mux_scbd_57.packet_count,57);
      packet_count_check(port_count[58],env.pf_vf_mux_scbd_58.packet_count,58);
      packet_count_check(port_count[59],env.pf_vf_mux_scbd_59.packet_count,59);
      packet_count_check(port_count[60],env.pf_vf_mux_scbd_60.packet_count,60);
      packet_count_check(port_count[61],env.pf_vf_mux_scbd_61.packet_count,61);
      packet_count_check(port_count[62],env.pf_vf_mux_scbd_62.packet_count,62);
      packet_count_check(port_count[63],env.pf_vf_mux_scbd_63.packet_count,63);
      packet_count_check(port_count[64],env.pf_vf_mux_scbd_64.packet_count,64);
      packet_count_check(port_count[65],env.pf_vf_mux_scbd_65.packet_count,65);
      packet_count_check(port_count[66],env.pf_vf_mux_scbd_66.packet_count,66);
      packet_count_check(port_count[67],env.pf_vf_mux_scbd_67.packet_count,67);
      packet_count_check(port_count[68],env.pf_vf_mux_scbd_68.packet_count,68);
      packet_count_check(port_count[69],env.pf_vf_mux_scbd_69.packet_count,69);
      packet_count_check(port_count[70],env.pf_vf_mux_scbd_70.packet_count,70);
      packet_count_check(port_count[71],env.pf_vf_mux_scbd_71.packet_count,71);
      packet_count_check(port_count[72],env.pf_vf_mux_scbd_72.packet_count,72);
      packet_count_check(port_count[73],env.pf_vf_mux_scbd_73.packet_count,73);
      packet_count_check(port_count[74],env.pf_vf_mux_scbd_74.packet_count,74);
      packet_count_check(port_count[75],env.pf_vf_mux_scbd_75.packet_count,75);
      packet_count_check(port_count[76],env.pf_vf_mux_scbd_76.packet_count,76);
      packet_count_check(port_count[77],env.pf_vf_mux_scbd_77.packet_count,77);
      packet_count_check(port_count[78],env.pf_vf_mux_scbd_78.packet_count,78);
      packet_count_check(port_count[79],env.pf_vf_mux_scbd_79.packet_count,79);
      packet_count_check(port_count[80],env.pf_vf_mux_scbd_80.packet_count,80);
      packet_count_check(port_count[81],env.pf_vf_mux_scbd_81.packet_count,81);
      packet_count_check(port_count[82],env.pf_vf_mux_scbd_82.packet_count,82);
      packet_count_check(port_count[83],env.pf_vf_mux_scbd_83.packet_count,83);
      packet_count_check(port_count[84],env.pf_vf_mux_scbd_84.packet_count,84);
      packet_count_check(port_count[85],env.pf_vf_mux_scbd_85.packet_count,85);
      packet_count_check(port_count[86],env.pf_vf_mux_scbd_86.packet_count,86);
      packet_count_check(port_count[87],env.pf_vf_mux_scbd_87.packet_count,87);
      packet_count_check(port_count[88],env.pf_vf_mux_scbd_88.packet_count,88);
      packet_count_check(port_count[89],env.pf_vf_mux_scbd_89.packet_count,89);
      packet_count_check(port_count[90],env.pf_vf_mux_scbd_90.packet_count,90);
      packet_count_check(port_count[91],env.pf_vf_mux_scbd_91.packet_count,91);
      packet_count_check(port_count[92],env.pf_vf_mux_scbd_92.packet_count,92);
      packet_count_check(port_count[93],env.pf_vf_mux_scbd_93.packet_count,93);
      packet_count_check(port_count[94],env.pf_vf_mux_scbd_94.packet_count,94);
      packet_count_check(port_count[95],env.pf_vf_mux_scbd_95.packet_count,95);
      packet_count_check(port_count[96],env.pf_vf_mux_scbd_96.packet_count,96);
      packet_count_check(port_count[97],env.pf_vf_mux_scbd_97.packet_count,97);
      packet_count_check(port_count[98],env.pf_vf_mux_scbd_98.packet_count,98);
      packet_count_check(port_count[99],env.pf_vf_mux_scbd_99.packet_count,99);
      packet_count_check(port_count[100],env.pf_vf_mux_scbd_100.packet_count,100);
      packet_count_check(port_count[101],env.pf_vf_mux_scbd_101.packet_count,101);
      packet_count_check(port_count[102],env.pf_vf_mux_scbd_102.packet_count,102);
      packet_count_check(port_count[103],env.pf_vf_mux_scbd_103.packet_count,103);
      packet_count_check(port_count[104],env.pf_vf_mux_scbd_104.packet_count,104);
      packet_count_check(port_count[105],env.pf_vf_mux_scbd_105.packet_count,105);
      packet_count_check(port_count[106],env.pf_vf_mux_scbd_106.packet_count,106);
      packet_count_check(port_count[107],env.pf_vf_mux_scbd_107.packet_count,107);
      packet_count_check(port_count[108],env.pf_vf_mux_scbd_108.packet_count,108);
      packet_count_check(port_count[109],env.pf_vf_mux_scbd_109.packet_count,109);
      packet_count_check(port_count[110],env.pf_vf_mux_scbd_110.packet_count,110);
      packet_count_check(port_count[111],env.pf_vf_mux_scbd_111.packet_count,111);
      packet_count_check(port_count[112],env.pf_vf_mux_scbd_112.packet_count,112);
      packet_count_check(port_count[113],env.pf_vf_mux_scbd_113.packet_count,113);
      packet_count_check(port_count[114],env.pf_vf_mux_scbd_114.packet_count,114);
      packet_count_check(port_count[115],env.pf_vf_mux_scbd_115.packet_count,115);
      packet_count_check(port_count[116],env.pf_vf_mux_scbd_116.packet_count,116);
      packet_count_check(port_count[117],env.pf_vf_mux_scbd_117.packet_count,117);
      packet_count_check(port_count[118],env.pf_vf_mux_scbd_118.packet_count,118);
      packet_count_check(port_count[119],env.pf_vf_mux_scbd_119.packet_count,119);
      packet_count_check(port_count[120],env.pf_vf_mux_scbd_120.packet_count,120);
      packet_count_check(port_count[121],env.pf_vf_mux_scbd_121.packet_count,121);
      packet_count_check(port_count[122],env.pf_vf_mux_scbd_122.packet_count,122);
      packet_count_check(port_count[123],env.pf_vf_mux_scbd_123.packet_count,123);
      packet_count_check(port_count[124],env.pf_vf_mux_scbd_124.packet_count,124);
      packet_count_check(port_count[125],env.pf_vf_mux_scbd_125.packet_count,125);
      packet_count_check(port_count[126],env.pf_vf_mux_scbd_126.packet_count,126);
      packet_count_check(port_count[127],env.pf_vf_mux_scbd_127.packet_count,127);
      packet_count_check(port_count[128],env.pf_vf_mux_scbd_128.packet_count,128);
      packet_count_check(port_count[129],env.pf_vf_mux_scbd_129.packet_count,129);
      packet_count_check(port_count[130],env.pf_vf_mux_scbd_130.packet_count,130);
      packet_count_check(port_count[131],env.pf_vf_mux_scbd_131.packet_count,131);
      packet_count_check(port_count[132],env.pf_vf_mux_scbd_132.packet_count,132);
      packet_count_check(port_count[133],env.pf_vf_mux_scbd_133.packet_count,133);
      packet_count_check(port_count[134],env.pf_vf_mux_scbd_134.packet_count,134);
      packet_count_check(port_count[135],env.pf_vf_mux_scbd_135.packet_count,135);
      packet_count_check(port_count[136],env.pf_vf_mux_scbd_136.packet_count,136);
      packet_count_check(port_count[137],env.pf_vf_mux_scbd_137.packet_count,137);
      packet_count_check(port_count[138],env.pf_vf_mux_scbd_138.packet_count,138);
      packet_count_check(port_count[139],env.pf_vf_mux_scbd_139.packet_count,139);
      packet_count_check(port_count[140],env.pf_vf_mux_scbd_140.packet_count,140);
      packet_count_check(port_count[141],env.pf_vf_mux_scbd_141.packet_count,141);
      packet_count_check(port_count[142],env.pf_vf_mux_scbd_142.packet_count,142);
      packet_count_check(port_count[143],env.pf_vf_mux_scbd_143.packet_count,143);
      packet_count_check(port_count[144],env.pf_vf_mux_scbd_144.packet_count,144);
      packet_count_check(port_count[145],env.pf_vf_mux_scbd_145.packet_count,145);
      packet_count_check(port_count[146],env.pf_vf_mux_scbd_146.packet_count,146);
      packet_count_check(port_count[147],env.pf_vf_mux_scbd_147.packet_count,147);
      packet_count_check(port_count[148],env.pf_vf_mux_scbd_148.packet_count,148);
      packet_count_check(port_count[149],env.pf_vf_mux_scbd_149.packet_count,149);
      packet_count_check(port_count[150],env.pf_vf_mux_scbd_150.packet_count,150);
      packet_count_check(port_count[151],env.pf_vf_mux_scbd_151.packet_count,151);
      packet_count_check(port_count[152],env.pf_vf_mux_scbd_152.packet_count,152);
      packet_count_check(port_count[153],env.pf_vf_mux_scbd_153.packet_count,153);
      packet_count_check(port_count[154],env.pf_vf_mux_scbd_154.packet_count,154);
      packet_count_check(port_count[155],env.pf_vf_mux_scbd_155.packet_count,155);
      packet_count_check(port_count[156],env.pf_vf_mux_scbd_156.packet_count,156);
      packet_count_check(port_count[157],env.pf_vf_mux_scbd_157.packet_count,157);
      packet_count_check(port_count[158],env.pf_vf_mux_scbd_158.packet_count,158);
      packet_count_check(port_count[159],env.pf_vf_mux_scbd_159.packet_count,159);
      packet_count_check(port_count[160],env.pf_vf_mux_scbd_160.packet_count,160);
      packet_count_check(port_count[161],env.pf_vf_mux_scbd_161.packet_count,161);
      packet_count_check(port_count[162],env.pf_vf_mux_scbd_162.packet_count,162);
      packet_count_check(port_count[163],env.pf_vf_mux_scbd_163.packet_count,163);
      packet_count_check(port_count[164],env.pf_vf_mux_scbd_164.packet_count,164);
      packet_count_check(port_count[165],env.pf_vf_mux_scbd_165.packet_count,165);
      packet_count_check(port_count[166],env.pf_vf_mux_scbd_166.packet_count,166);
      packet_count_check(port_count[167],env.pf_vf_mux_scbd_167.packet_count,167);
      packet_count_check(port_count[168],env.pf_vf_mux_scbd_168.packet_count,168);
      packet_count_check(port_count[169],env.pf_vf_mux_scbd_169.packet_count,169);
      packet_count_check(port_count[170],env.pf_vf_mux_scbd_170.packet_count,170);
      packet_count_check(port_count[171],env.pf_vf_mux_scbd_171.packet_count,171);
      packet_count_check(port_count[172],env.pf_vf_mux_scbd_172.packet_count,172);
      packet_count_check(port_count[173],env.pf_vf_mux_scbd_173.packet_count,173);
      packet_count_check(port_count[174],env.pf_vf_mux_scbd_174.packet_count,174);
      packet_count_check(port_count[175],env.pf_vf_mux_scbd_175.packet_count,175);
      packet_count_check(port_count[176],env.pf_vf_mux_scbd_176.packet_count,176);
      packet_count_check(port_count[177],env.pf_vf_mux_scbd_177.packet_count,177);
      packet_count_check(port_count[178],env.pf_vf_mux_scbd_178.packet_count,178);
      packet_count_check(port_count[179],env.pf_vf_mux_scbd_179.packet_count,179);
      packet_count_check(port_count[180],env.pf_vf_mux_scbd_180.packet_count,180);
      packet_count_check(port_count[181],env.pf_vf_mux_scbd_181.packet_count,181);
      packet_count_check(port_count[182],env.pf_vf_mux_scbd_182.packet_count,182);
      packet_count_check(port_count[183],env.pf_vf_mux_scbd_183.packet_count,183);
      packet_count_check(port_count[184],env.pf_vf_mux_scbd_184.packet_count,184);
      packet_count_check(port_count[185],env.pf_vf_mux_scbd_185.packet_count,185);
      packet_count_check(port_count[186],env.pf_vf_mux_scbd_186.packet_count,186);
      packet_count_check(port_count[187],env.pf_vf_mux_scbd_187.packet_count,187);
      packet_count_check(port_count[188],env.pf_vf_mux_scbd_188.packet_count,188);
      packet_count_check(port_count[189],env.pf_vf_mux_scbd_189.packet_count,189);
      packet_count_check(port_count[190],env.pf_vf_mux_scbd_190.packet_count,190);
      packet_count_check(port_count[191],env.pf_vf_mux_scbd_191.packet_count,191);
      packet_count_check(port_count[192],env.pf_vf_mux_scbd_192.packet_count,192);
      packet_count_check(port_count[193],env.pf_vf_mux_scbd_193.packet_count,193);
      packet_count_check(port_count[194],env.pf_vf_mux_scbd_194.packet_count,194);
      packet_count_check(port_count[195],env.pf_vf_mux_scbd_195.packet_count,195);
      packet_count_check(port_count[196],env.pf_vf_mux_scbd_196.packet_count,196);
      packet_count_check(port_count[197],env.pf_vf_mux_scbd_197.packet_count,197);
      packet_count_check(port_count[198],env.pf_vf_mux_scbd_198.packet_count,198);
      packet_count_check(port_count[199],env.pf_vf_mux_scbd_199.packet_count,199);
      packet_count_check(port_count[200],env.pf_vf_mux_scbd_200.packet_count,200);
      packet_count_check(port_count[201],env.pf_vf_mux_scbd_201.packet_count,201);
      packet_count_check(port_count[202],env.pf_vf_mux_scbd_202.packet_count,202);
      packet_count_check(port_count[203],env.pf_vf_mux_scbd_203.packet_count,203);
      packet_count_check(port_count[204],env.pf_vf_mux_scbd_204.packet_count,204);
      packet_count_check(port_count[205],env.pf_vf_mux_scbd_205.packet_count,205);
      packet_count_check(port_count[206],env.pf_vf_mux_scbd_206.packet_count,206);
      packet_count_check(port_count[207],env.pf_vf_mux_scbd_207.packet_count,207);
      packet_count_check(port_count[208],env.pf_vf_mux_scbd_208.packet_count,208);
      packet_count_check(port_count[209],env.pf_vf_mux_scbd_209.packet_count,209);
      packet_count_check(port_count[210],env.pf_vf_mux_scbd_210.packet_count,210);
      packet_count_check(port_count[211],env.pf_vf_mux_scbd_211.packet_count,211);
      packet_count_check(port_count[212],env.pf_vf_mux_scbd_212.packet_count,212);
      packet_count_check(port_count[213],env.pf_vf_mux_scbd_213.packet_count,213);
      packet_count_check(port_count[214],env.pf_vf_mux_scbd_214.packet_count,214);
      packet_count_check(port_count[215],env.pf_vf_mux_scbd_215.packet_count,215);
      packet_count_check(port_count[216],env.pf_vf_mux_scbd_216.packet_count,216);
      packet_count_check(port_count[217],env.pf_vf_mux_scbd_217.packet_count,217);
      packet_count_check(port_count[218],env.pf_vf_mux_scbd_218.packet_count,218);
      packet_count_check(port_count[219],env.pf_vf_mux_scbd_219.packet_count,219);
      packet_count_check(port_count[220],env.pf_vf_mux_scbd_220.packet_count,220);
      packet_count_check(port_count[221],env.pf_vf_mux_scbd_221.packet_count,221);
      packet_count_check(port_count[222],env.pf_vf_mux_scbd_222.packet_count,222);
      packet_count_check(port_count[223],env.pf_vf_mux_scbd_223.packet_count,223);
      packet_count_check(port_count[224],env.pf_vf_mux_scbd_224.packet_count,224);
      packet_count_check(port_count[225],env.pf_vf_mux_scbd_225.packet_count,225);
      packet_count_check(port_count[226],env.pf_vf_mux_scbd_226.packet_count,226);
      packet_count_check(port_count[227],env.pf_vf_mux_scbd_227.packet_count,227);
      packet_count_check(port_count[228],env.pf_vf_mux_scbd_228.packet_count,228);
      packet_count_check(port_count[229],env.pf_vf_mux_scbd_229.packet_count,229);
      packet_count_check(port_count[230],env.pf_vf_mux_scbd_230.packet_count,230);
      packet_count_check(port_count[231],env.pf_vf_mux_scbd_231.packet_count,231);
      packet_count_check(port_count[232],env.pf_vf_mux_scbd_232.packet_count,232);
      packet_count_check(port_count[233],env.pf_vf_mux_scbd_233.packet_count,233);
      packet_count_check(port_count[234],env.pf_vf_mux_scbd_234.packet_count,234);
      packet_count_check(port_count[235],env.pf_vf_mux_scbd_235.packet_count,235);
      packet_count_check(port_count[236],env.pf_vf_mux_scbd_236.packet_count,236);
      packet_count_check(port_count[237],env.pf_vf_mux_scbd_237.packet_count,237);
      packet_count_check(port_count[238],env.pf_vf_mux_scbd_238.packet_count,238);
      packet_count_check(port_count[239],env.pf_vf_mux_scbd_239.packet_count,239);
      packet_count_check(port_count[240],env.pf_vf_mux_scbd_240.packet_count,240);
      packet_count_check(port_count[241],env.pf_vf_mux_scbd_241.packet_count,241);
      packet_count_check(port_count[242],env.pf_vf_mux_scbd_242.packet_count,242);
      packet_count_check(port_count[243],env.pf_vf_mux_scbd_243.packet_count,243);
      packet_count_check(port_count[244],env.pf_vf_mux_scbd_244.packet_count,244);
      packet_count_check(port_count[245],env.pf_vf_mux_scbd_245.packet_count,245);
      packet_count_check(port_count[246],env.pf_vf_mux_scbd_246.packet_count,246);
      packet_count_check(port_count[247],env.pf_vf_mux_scbd_247.packet_count,247);
      packet_count_check(port_count[248],env.pf_vf_mux_scbd_248.packet_count,248);
      packet_count_check(port_count[249],env.pf_vf_mux_scbd_249.packet_count,249);
      packet_count_check(port_count[250],env.pf_vf_mux_scbd_250.packet_count,250);
      packet_count_check(port_count[251],env.pf_vf_mux_scbd_251.packet_count,251);
      packet_count_check(port_count[252],env.pf_vf_mux_scbd_252.packet_count,252);
      packet_count_check(port_count[253],env.pf_vf_mux_scbd_253.packet_count,253);
      packet_count_check(port_count[254],env.pf_vf_mux_scbd_254.packet_count,254);
      packet_count_check(port_count[255],env.pf_vf_mux_scbd_255.packet_count,255);
      packet_count_check(port_count[256],env.pf_vf_mux_scbd_256.packet_count,256);
      packet_count_check(port_count[257],env.pf_vf_mux_scbd_257.packet_count,257);
      packet_count_check(port_count[258],env.pf_vf_mux_scbd_258.packet_count,258);
      packet_count_check(port_count[259],env.pf_vf_mux_scbd_259.packet_count,259);
      packet_count_check(port_count[260],env.pf_vf_mux_scbd_260.packet_count,260);
      packet_count_check(port_count[261],env.pf_vf_mux_scbd_261.packet_count,261);
      packet_count_check(port_count[262],env.pf_vf_mux_scbd_262.packet_count,262);
      packet_count_check(port_count[263],env.pf_vf_mux_scbd_263.packet_count,263);
      packet_count_check(port_count[264],env.pf_vf_mux_scbd_264.packet_count,264);
      packet_count_check(port_count[265],env.pf_vf_mux_scbd_265.packet_count,265);
      packet_count_check(port_count[266],env.pf_vf_mux_scbd_266.packet_count,266);
      packet_count_check(port_count[267],env.pf_vf_mux_scbd_267.packet_count,267);
      packet_count_check(port_count[268],env.pf_vf_mux_scbd_268.packet_count,268);
      packet_count_check(port_count[269],env.pf_vf_mux_scbd_269.packet_count,269);
      packet_count_check(port_count[270],env.pf_vf_mux_scbd_270.packet_count,270);
      packet_count_check(port_count[271],env.pf_vf_mux_scbd_271.packet_count,271);
      packet_count_check(port_count[272],env.pf_vf_mux_scbd_272.packet_count,272);
      packet_count_check(port_count[273],env.pf_vf_mux_scbd_273.packet_count,273);
      packet_count_check(port_count[274],env.pf_vf_mux_scbd_274.packet_count,274);
      packet_count_check(port_count[275],env.pf_vf_mux_scbd_275.packet_count,275);
      packet_count_check(port_count[276],env.pf_vf_mux_scbd_276.packet_count,276);
      packet_count_check(port_count[277],env.pf_vf_mux_scbd_277.packet_count,277);
      packet_count_check(port_count[278],env.pf_vf_mux_scbd_278.packet_count,278);
      packet_count_check(port_count[279],env.pf_vf_mux_scbd_279.packet_count,279);
      packet_count_check(port_count[280],env.pf_vf_mux_scbd_280.packet_count,280);
      packet_count_check(port_count[281],env.pf_vf_mux_scbd_281.packet_count,281);
      packet_count_check(port_count[282],env.pf_vf_mux_scbd_282.packet_count,282);
      packet_count_check(port_count[283],env.pf_vf_mux_scbd_283.packet_count,283);
      packet_count_check(port_count[284],env.pf_vf_mux_scbd_284.packet_count,284);
      packet_count_check(port_count[285],env.pf_vf_mux_scbd_285.packet_count,285);
      packet_count_check(port_count[286],env.pf_vf_mux_scbd_286.packet_count,286);
      packet_count_check(port_count[287],env.pf_vf_mux_scbd_287.packet_count,287);
      packet_count_check(port_count[288],env.pf_vf_mux_scbd_288.packet_count,288);
      packet_count_check(port_count[289],env.pf_vf_mux_scbd_289.packet_count,289);
      packet_count_check(port_count[290],env.pf_vf_mux_scbd_290.packet_count,290);
      packet_count_check(port_count[291],env.pf_vf_mux_scbd_291.packet_count,291);
      packet_count_check(port_count[292],env.pf_vf_mux_scbd_292.packet_count,292);
      packet_count_check(port_count[293],env.pf_vf_mux_scbd_293.packet_count,293);
      packet_count_check(port_count[294],env.pf_vf_mux_scbd_294.packet_count,294);
      packet_count_check(port_count[295],env.pf_vf_mux_scbd_295.packet_count,295);
      packet_count_check(port_count[296],env.pf_vf_mux_scbd_296.packet_count,296);
      packet_count_check(port_count[297],env.pf_vf_mux_scbd_297.packet_count,297);
      packet_count_check(port_count[298],env.pf_vf_mux_scbd_298.packet_count,298);
      packet_count_check(port_count[299],env.pf_vf_mux_scbd_299.packet_count,299);
      packet_count_check(port_count[300],env.pf_vf_mux_scbd_300.packet_count,300);
      packet_count_check(port_count[301],env.pf_vf_mux_scbd_301.packet_count,301);
      packet_count_check(port_count[302],env.pf_vf_mux_scbd_302.packet_count,302);
      packet_count_check(port_count[303],env.pf_vf_mux_scbd_303.packet_count,303);
      packet_count_check(port_count[304],env.pf_vf_mux_scbd_304.packet_count,304);
      packet_count_check(port_count[305],env.pf_vf_mux_scbd_305.packet_count,305);
      packet_count_check(port_count[306],env.pf_vf_mux_scbd_306.packet_count,306);
      packet_count_check(port_count[307],env.pf_vf_mux_scbd_307.packet_count,307);
      packet_count_check(port_count[308],env.pf_vf_mux_scbd_308.packet_count,308);
      packet_count_check(port_count[309],env.pf_vf_mux_scbd_309.packet_count,309);
      packet_count_check(port_count[310],env.pf_vf_mux_scbd_310.packet_count,310);
      packet_count_check(port_count[311],env.pf_vf_mux_scbd_311.packet_count,311);
      packet_count_check(port_count[312],env.pf_vf_mux_scbd_312.packet_count,312);
      packet_count_check(port_count[313],env.pf_vf_mux_scbd_313.packet_count,313);
      packet_count_check(port_count[314],env.pf_vf_mux_scbd_314.packet_count,314);
      packet_count_check(port_count[315],env.pf_vf_mux_scbd_315.packet_count,315);
      packet_count_check(port_count[316],env.pf_vf_mux_scbd_316.packet_count,316);
      packet_count_check(port_count[317],env.pf_vf_mux_scbd_317.packet_count,317);
      packet_count_check(port_count[318],env.pf_vf_mux_scbd_318.packet_count,318);
      packet_count_check(port_count[319],env.pf_vf_mux_scbd_319.packet_count,319);
      packet_count_check(port_count[320],env.pf_vf_mux_scbd_320.packet_count,320);
      packet_count_check(port_count[321],env.pf_vf_mux_scbd_321.packet_count,321);
      packet_count_check(port_count[322],env.pf_vf_mux_scbd_322.packet_count,322);
      packet_count_check(port_count[323],env.pf_vf_mux_scbd_323.packet_count,323);
      packet_count_check(port_count[324],env.pf_vf_mux_scbd_324.packet_count,324);
      packet_count_check(port_count[325],env.pf_vf_mux_scbd_325.packet_count,325);
      packet_count_check(port_count[326],env.pf_vf_mux_scbd_326.packet_count,326);
      packet_count_check(port_count[327],env.pf_vf_mux_scbd_327.packet_count,327);
      packet_count_check(port_count[328],env.pf_vf_mux_scbd_328.packet_count,328);
      packet_count_check(port_count[329],env.pf_vf_mux_scbd_329.packet_count,329);
      packet_count_check(port_count[330],env.pf_vf_mux_scbd_330.packet_count,330);
      packet_count_check(port_count[331],env.pf_vf_mux_scbd_331.packet_count,331);
      packet_count_check(port_count[332],env.pf_vf_mux_scbd_332.packet_count,332);
      packet_count_check(port_count[333],env.pf_vf_mux_scbd_333.packet_count,333);
      packet_count_check(port_count[334],env.pf_vf_mux_scbd_334.packet_count,334);
      packet_count_check(port_count[335],env.pf_vf_mux_scbd_335.packet_count,335);
      packet_count_check(port_count[336],env.pf_vf_mux_scbd_336.packet_count,336);
      packet_count_check(port_count[337],env.pf_vf_mux_scbd_337.packet_count,337);
      packet_count_check(port_count[338],env.pf_vf_mux_scbd_338.packet_count,338);
      packet_count_check(port_count[339],env.pf_vf_mux_scbd_339.packet_count,339);
      packet_count_check(port_count[340],env.pf_vf_mux_scbd_340.packet_count,340);
      packet_count_check(port_count[341],env.pf_vf_mux_scbd_341.packet_count,341);
      packet_count_check(port_count[342],env.pf_vf_mux_scbd_342.packet_count,342);
      packet_count_check(port_count[343],env.pf_vf_mux_scbd_343.packet_count,343);
      packet_count_check(port_count[344],env.pf_vf_mux_scbd_344.packet_count,344);
      packet_count_check(port_count[345],env.pf_vf_mux_scbd_345.packet_count,345);
      packet_count_check(port_count[346],env.pf_vf_mux_scbd_346.packet_count,346);
      packet_count_check(port_count[347],env.pf_vf_mux_scbd_347.packet_count,347);
      packet_count_check(port_count[348],env.pf_vf_mux_scbd_348.packet_count,348);
      packet_count_check(port_count[349],env.pf_vf_mux_scbd_349.packet_count,349);
      packet_count_check(port_count[350],env.pf_vf_mux_scbd_350.packet_count,350);
      packet_count_check(port_count[351],env.pf_vf_mux_scbd_351.packet_count,351);
      packet_count_check(port_count[352],env.pf_vf_mux_scbd_352.packet_count,352);
      packet_count_check(port_count[353],env.pf_vf_mux_scbd_353.packet_count,353);
      packet_count_check(port_count[354],env.pf_vf_mux_scbd_354.packet_count,354);
      packet_count_check(port_count[355],env.pf_vf_mux_scbd_355.packet_count,355);
      packet_count_check(port_count[356],env.pf_vf_mux_scbd_356.packet_count,356);
      packet_count_check(port_count[357],env.pf_vf_mux_scbd_357.packet_count,357);
      packet_count_check(port_count[358],env.pf_vf_mux_scbd_358.packet_count,358);
      packet_count_check(port_count[359],env.pf_vf_mux_scbd_359.packet_count,359);
      packet_count_check(port_count[360],env.pf_vf_mux_scbd_360.packet_count,360);
      packet_count_check(port_count[361],env.pf_vf_mux_scbd_361.packet_count,361);
      packet_count_check(port_count[362],env.pf_vf_mux_scbd_362.packet_count,362);
      packet_count_check(port_count[363],env.pf_vf_mux_scbd_363.packet_count,363);
      packet_count_check(port_count[364],env.pf_vf_mux_scbd_364.packet_count,364);
      packet_count_check(port_count[365],env.pf_vf_mux_scbd_365.packet_count,365);
      packet_count_check(port_count[366],env.pf_vf_mux_scbd_366.packet_count,366);
      packet_count_check(port_count[367],env.pf_vf_mux_scbd_367.packet_count,367);
      packet_count_check(port_count[368],env.pf_vf_mux_scbd_368.packet_count,368);
      packet_count_check(port_count[369],env.pf_vf_mux_scbd_369.packet_count,369);
      packet_count_check(port_count[370],env.pf_vf_mux_scbd_370.packet_count,370);
      packet_count_check(port_count[371],env.pf_vf_mux_scbd_371.packet_count,371);
      packet_count_check(port_count[372],env.pf_vf_mux_scbd_372.packet_count,372);
      packet_count_check(port_count[373],env.pf_vf_mux_scbd_373.packet_count,373);
      packet_count_check(port_count[374],env.pf_vf_mux_scbd_374.packet_count,374);
      packet_count_check(port_count[375],env.pf_vf_mux_scbd_375.packet_count,375);
      packet_count_check(port_count[376],env.pf_vf_mux_scbd_376.packet_count,376);
      packet_count_check(port_count[377],env.pf_vf_mux_scbd_377.packet_count,377);
      packet_count_check(port_count[378],env.pf_vf_mux_scbd_378.packet_count,378);
      packet_count_check(port_count[379],env.pf_vf_mux_scbd_379.packet_count,379);
      packet_count_check(port_count[380],env.pf_vf_mux_scbd_380.packet_count,380);
      packet_count_check(port_count[381],env.pf_vf_mux_scbd_381.packet_count,381);
      packet_count_check(port_count[382],env.pf_vf_mux_scbd_382.packet_count,382);
      packet_count_check(port_count[383],env.pf_vf_mux_scbd_383.packet_count,383);
      packet_count_check(port_count[384],env.pf_vf_mux_scbd_384.packet_count,384);
      packet_count_check(port_count[385],env.pf_vf_mux_scbd_385.packet_count,385);
      packet_count_check(port_count[386],env.pf_vf_mux_scbd_386.packet_count,386);
      packet_count_check(port_count[387],env.pf_vf_mux_scbd_387.packet_count,387);
      packet_count_check(port_count[388],env.pf_vf_mux_scbd_388.packet_count,388);
      packet_count_check(port_count[389],env.pf_vf_mux_scbd_389.packet_count,389);
      packet_count_check(port_count[390],env.pf_vf_mux_scbd_390.packet_count,390);
      packet_count_check(port_count[391],env.pf_vf_mux_scbd_391.packet_count,391);
      packet_count_check(port_count[392],env.pf_vf_mux_scbd_392.packet_count,392);
      packet_count_check(port_count[393],env.pf_vf_mux_scbd_393.packet_count,393);
      packet_count_check(port_count[394],env.pf_vf_mux_scbd_394.packet_count,394);
      packet_count_check(port_count[395],env.pf_vf_mux_scbd_395.packet_count,395);
      packet_count_check(port_count[396],env.pf_vf_mux_scbd_396.packet_count,396);
      packet_count_check(port_count[397],env.pf_vf_mux_scbd_397.packet_count,397);
      packet_count_check(port_count[398],env.pf_vf_mux_scbd_398.packet_count,398);
      packet_count_check(port_count[399],env.pf_vf_mux_scbd_399.packet_count,399);
      packet_count_check(port_count[400],env.pf_vf_mux_scbd_400.packet_count,400);
      packet_count_check(port_count[401],env.pf_vf_mux_scbd_401.packet_count,401);
      packet_count_check(port_count[402],env.pf_vf_mux_scbd_402.packet_count,402);
      packet_count_check(port_count[403],env.pf_vf_mux_scbd_403.packet_count,403);
      packet_count_check(port_count[404],env.pf_vf_mux_scbd_404.packet_count,404);
      packet_count_check(port_count[405],env.pf_vf_mux_scbd_405.packet_count,405);
      packet_count_check(port_count[406],env.pf_vf_mux_scbd_406.packet_count,406);
      packet_count_check(port_count[407],env.pf_vf_mux_scbd_407.packet_count,407);
      packet_count_check(port_count[408],env.pf_vf_mux_scbd_408.packet_count,408);
      packet_count_check(port_count[409],env.pf_vf_mux_scbd_409.packet_count,409);
      packet_count_check(port_count[410],env.pf_vf_mux_scbd_410.packet_count,410);
      packet_count_check(port_count[411],env.pf_vf_mux_scbd_411.packet_count,411);
      packet_count_check(port_count[412],env.pf_vf_mux_scbd_412.packet_count,412);
      packet_count_check(port_count[413],env.pf_vf_mux_scbd_413.packet_count,413);
      packet_count_check(port_count[414],env.pf_vf_mux_scbd_414.packet_count,414);
      packet_count_check(port_count[415],env.pf_vf_mux_scbd_415.packet_count,415);
      packet_count_check(port_count[416],env.pf_vf_mux_scbd_416.packet_count,416);
      packet_count_check(port_count[417],env.pf_vf_mux_scbd_417.packet_count,417);
      packet_count_check(port_count[418],env.pf_vf_mux_scbd_418.packet_count,418);
      packet_count_check(port_count[419],env.pf_vf_mux_scbd_419.packet_count,419);
      packet_count_check(port_count[420],env.pf_vf_mux_scbd_420.packet_count,420);
      packet_count_check(port_count[421],env.pf_vf_mux_scbd_421.packet_count,421);
      packet_count_check(port_count[422],env.pf_vf_mux_scbd_422.packet_count,422);
      packet_count_check(port_count[423],env.pf_vf_mux_scbd_423.packet_count,423);
      packet_count_check(port_count[424],env.pf_vf_mux_scbd_424.packet_count,424);
      packet_count_check(port_count[425],env.pf_vf_mux_scbd_425.packet_count,425);
      packet_count_check(port_count[426],env.pf_vf_mux_scbd_426.packet_count,426);
      packet_count_check(port_count[427],env.pf_vf_mux_scbd_427.packet_count,427);
      packet_count_check(port_count[428],env.pf_vf_mux_scbd_428.packet_count,428);
      packet_count_check(port_count[429],env.pf_vf_mux_scbd_429.packet_count,429);
      packet_count_check(port_count[430],env.pf_vf_mux_scbd_430.packet_count,430);
      packet_count_check(port_count[431],env.pf_vf_mux_scbd_431.packet_count,431);
      packet_count_check(port_count[432],env.pf_vf_mux_scbd_432.packet_count,432);
      packet_count_check(port_count[433],env.pf_vf_mux_scbd_433.packet_count,433);
      packet_count_check(port_count[434],env.pf_vf_mux_scbd_434.packet_count,434);
      packet_count_check(port_count[435],env.pf_vf_mux_scbd_435.packet_count,435);
      packet_count_check(port_count[436],env.pf_vf_mux_scbd_436.packet_count,436);
      packet_count_check(port_count[437],env.pf_vf_mux_scbd_437.packet_count,437);
      packet_count_check(port_count[438],env.pf_vf_mux_scbd_438.packet_count,438);
      packet_count_check(port_count[439],env.pf_vf_mux_scbd_439.packet_count,439);
      packet_count_check(port_count[440],env.pf_vf_mux_scbd_440.packet_count,440);
      packet_count_check(port_count[441],env.pf_vf_mux_scbd_441.packet_count,441);
      packet_count_check(port_count[442],env.pf_vf_mux_scbd_442.packet_count,442);
      packet_count_check(port_count[443],env.pf_vf_mux_scbd_443.packet_count,443);
      packet_count_check(port_count[444],env.pf_vf_mux_scbd_444.packet_count,444);
      packet_count_check(port_count[445],env.pf_vf_mux_scbd_445.packet_count,445);
      packet_count_check(port_count[446],env.pf_vf_mux_scbd_446.packet_count,446);
      packet_count_check(port_count[447],env.pf_vf_mux_scbd_447.packet_count,447);
      packet_count_check(port_count[448],env.pf_vf_mux_scbd_448.packet_count,448);
      packet_count_check(port_count[449],env.pf_vf_mux_scbd_449.packet_count,449);
      packet_count_check(port_count[450],env.pf_vf_mux_scbd_450.packet_count,450);
      packet_count_check(port_count[451],env.pf_vf_mux_scbd_451.packet_count,451);
      packet_count_check(port_count[452],env.pf_vf_mux_scbd_452.packet_count,452);
      packet_count_check(port_count[453],env.pf_vf_mux_scbd_453.packet_count,453);
      packet_count_check(port_count[454],env.pf_vf_mux_scbd_454.packet_count,454);
      packet_count_check(port_count[455],env.pf_vf_mux_scbd_455.packet_count,455);
      packet_count_check(port_count[456],env.pf_vf_mux_scbd_456.packet_count,456);
      packet_count_check(port_count[457],env.pf_vf_mux_scbd_457.packet_count,457);
      packet_count_check(port_count[458],env.pf_vf_mux_scbd_458.packet_count,458);
      packet_count_check(port_count[459],env.pf_vf_mux_scbd_459.packet_count,459);
      packet_count_check(port_count[460],env.pf_vf_mux_scbd_460.packet_count,460);
      packet_count_check(port_count[461],env.pf_vf_mux_scbd_461.packet_count,461);
      packet_count_check(port_count[462],env.pf_vf_mux_scbd_462.packet_count,462);
      packet_count_check(port_count[463],env.pf_vf_mux_scbd_463.packet_count,463);
      packet_count_check(port_count[464],env.pf_vf_mux_scbd_464.packet_count,464);
      packet_count_check(port_count[465],env.pf_vf_mux_scbd_465.packet_count,465);
      packet_count_check(port_count[466],env.pf_vf_mux_scbd_466.packet_count,466);
      packet_count_check(port_count[467],env.pf_vf_mux_scbd_467.packet_count,467);
      packet_count_check(port_count[468],env.pf_vf_mux_scbd_468.packet_count,468);
      packet_count_check(port_count[469],env.pf_vf_mux_scbd_469.packet_count,469);
      packet_count_check(port_count[470],env.pf_vf_mux_scbd_470.packet_count,470);
      packet_count_check(port_count[471],env.pf_vf_mux_scbd_471.packet_count,471);
      packet_count_check(port_count[472],env.pf_vf_mux_scbd_472.packet_count,472);
      packet_count_check(port_count[473],env.pf_vf_mux_scbd_473.packet_count,473);
      packet_count_check(port_count[474],env.pf_vf_mux_scbd_474.packet_count,474);
      packet_count_check(port_count[475],env.pf_vf_mux_scbd_475.packet_count,475);
      packet_count_check(port_count[476],env.pf_vf_mux_scbd_476.packet_count,476);
      packet_count_check(port_count[477],env.pf_vf_mux_scbd_477.packet_count,477);
      packet_count_check(port_count[478],env.pf_vf_mux_scbd_478.packet_count,478);
      packet_count_check(port_count[479],env.pf_vf_mux_scbd_479.packet_count,479);
      packet_count_check(port_count[480],env.pf_vf_mux_scbd_480.packet_count,480);
      packet_count_check(port_count[481],env.pf_vf_mux_scbd_481.packet_count,481);
      packet_count_check(port_count[482],env.pf_vf_mux_scbd_482.packet_count,482);
      packet_count_check(port_count[483],env.pf_vf_mux_scbd_483.packet_count,483);
      packet_count_check(port_count[484],env.pf_vf_mux_scbd_484.packet_count,484);
      packet_count_check(port_count[485],env.pf_vf_mux_scbd_485.packet_count,485);
      packet_count_check(port_count[486],env.pf_vf_mux_scbd_486.packet_count,486);
      packet_count_check(port_count[487],env.pf_vf_mux_scbd_487.packet_count,487);
      packet_count_check(port_count[488],env.pf_vf_mux_scbd_488.packet_count,488);
      packet_count_check(port_count[489],env.pf_vf_mux_scbd_489.packet_count,489);
      packet_count_check(port_count[490],env.pf_vf_mux_scbd_490.packet_count,490);
      packet_count_check(port_count[491],env.pf_vf_mux_scbd_491.packet_count,491);
      packet_count_check(port_count[492],env.pf_vf_mux_scbd_492.packet_count,492);
      packet_count_check(port_count[493],env.pf_vf_mux_scbd_493.packet_count,493);
      packet_count_check(port_count[494],env.pf_vf_mux_scbd_494.packet_count,494);
      packet_count_check(port_count[495],env.pf_vf_mux_scbd_495.packet_count,495);
      packet_count_check(port_count[496],env.pf_vf_mux_scbd_496.packet_count,496);
      packet_count_check(port_count[497],env.pf_vf_mux_scbd_497.packet_count,497);
      packet_count_check(port_count[498],env.pf_vf_mux_scbd_498.packet_count,498);
      packet_count_check(port_count[499],env.pf_vf_mux_scbd_499.packet_count,499);
      packet_count_check(port_count[500],env.pf_vf_mux_scbd_500.packet_count,500);
      packet_count_check(port_count[501],env.pf_vf_mux_scbd_501.packet_count,501);
      packet_count_check(port_count[502],env.pf_vf_mux_scbd_502.packet_count,502);
      packet_count_check(port_count[503],env.pf_vf_mux_scbd_503.packet_count,503);
      packet_count_check(port_count[504],env.pf_vf_mux_scbd_504.packet_count,504);
      packet_count_check(port_count[505],env.pf_vf_mux_scbd_505.packet_count,505);
      packet_count_check(port_count[506],env.pf_vf_mux_scbd_506.packet_count,506);
      packet_count_check(port_count[507],env.pf_vf_mux_scbd_507.packet_count,507);
      packet_count_check(port_count[508],env.pf_vf_mux_scbd_508.packet_count,508);
      packet_count_check(port_count[509],env.pf_vf_mux_scbd_509.packet_count,509);
      packet_count_check(port_count[510],env.pf_vf_mux_scbd_510.packet_count,510);
      packet_count_check(port_count[511],env.pf_vf_mux_scbd_511.packet_count,511);
      packet_count_check(port_count[512],env.pf_vf_mux_scbd_512.packet_count,512);
      packet_count_check(port_count[513],env.pf_vf_mux_scbd_513.packet_count,513);
      packet_count_check(port_count[514],env.pf_vf_mux_scbd_514.packet_count,514);
      packet_count_check(port_count[515],env.pf_vf_mux_scbd_515.packet_count,515);
      packet_count_check(port_count[516],env.pf_vf_mux_scbd_516.packet_count,516);
      packet_count_check(port_count[517],env.pf_vf_mux_scbd_517.packet_count,517);
      packet_count_check(port_count[518],env.pf_vf_mux_scbd_518.packet_count,518);
      packet_count_check(port_count[519],env.pf_vf_mux_scbd_519.packet_count,519);
      packet_count_check(port_count[520],env.pf_vf_mux_scbd_520.packet_count,520);
      packet_count_check(port_count[521],env.pf_vf_mux_scbd_521.packet_count,521);
      packet_count_check(port_count[522],env.pf_vf_mux_scbd_522.packet_count,522);
      packet_count_check(port_count[523],env.pf_vf_mux_scbd_523.packet_count,523);
      packet_count_check(port_count[524],env.pf_vf_mux_scbd_524.packet_count,524);
      packet_count_check(port_count[525],env.pf_vf_mux_scbd_525.packet_count,525);
      packet_count_check(port_count[526],env.pf_vf_mux_scbd_526.packet_count,526);
      packet_count_check(port_count[527],env.pf_vf_mux_scbd_527.packet_count,527);
      packet_count_check(port_count[528],env.pf_vf_mux_scbd_528.packet_count,528);
      packet_count_check(port_count[529],env.pf_vf_mux_scbd_529.packet_count,529);
      packet_count_check(port_count[530],env.pf_vf_mux_scbd_530.packet_count,530);
      packet_count_check(port_count[531],env.pf_vf_mux_scbd_531.packet_count,531);
      packet_count_check(port_count[532],env.pf_vf_mux_scbd_532.packet_count,532);
      packet_count_check(port_count[533],env.pf_vf_mux_scbd_533.packet_count,533);
      packet_count_check(port_count[534],env.pf_vf_mux_scbd_534.packet_count,534);
      packet_count_check(port_count[535],env.pf_vf_mux_scbd_535.packet_count,535);
      packet_count_check(port_count[536],env.pf_vf_mux_scbd_536.packet_count,536);
      packet_count_check(port_count[537],env.pf_vf_mux_scbd_537.packet_count,537);
      packet_count_check(port_count[538],env.pf_vf_mux_scbd_538.packet_count,538);
      packet_count_check(port_count[539],env.pf_vf_mux_scbd_539.packet_count,539);
      packet_count_check(port_count[540],env.pf_vf_mux_scbd_540.packet_count,540);
      packet_count_check(port_count[541],env.pf_vf_mux_scbd_541.packet_count,541);
      packet_count_check(port_count[542],env.pf_vf_mux_scbd_542.packet_count,542);
      packet_count_check(port_count[543],env.pf_vf_mux_scbd_543.packet_count,543);
      packet_count_check(port_count[544],env.pf_vf_mux_scbd_544.packet_count,544);
      packet_count_check(port_count[545],env.pf_vf_mux_scbd_545.packet_count,545);
      packet_count_check(port_count[546],env.pf_vf_mux_scbd_546.packet_count,546);
      packet_count_check(port_count[547],env.pf_vf_mux_scbd_547.packet_count,547);
      packet_count_check(port_count[548],env.pf_vf_mux_scbd_548.packet_count,548);
      packet_count_check(port_count[549],env.pf_vf_mux_scbd_549.packet_count,549);
      packet_count_check(port_count[550],env.pf_vf_mux_scbd_550.packet_count,550);
      packet_count_check(port_count[551],env.pf_vf_mux_scbd_551.packet_count,551);
      packet_count_check(port_count[552],env.pf_vf_mux_scbd_552.packet_count,552);
      packet_count_check(port_count[553],env.pf_vf_mux_scbd_553.packet_count,553);
      packet_count_check(port_count[554],env.pf_vf_mux_scbd_554.packet_count,554);
      packet_count_check(port_count[555],env.pf_vf_mux_scbd_555.packet_count,555);
      packet_count_check(port_count[556],env.pf_vf_mux_scbd_556.packet_count,556);
      packet_count_check(port_count[557],env.pf_vf_mux_scbd_557.packet_count,557);
      packet_count_check(port_count[558],env.pf_vf_mux_scbd_558.packet_count,558);
      packet_count_check(port_count[559],env.pf_vf_mux_scbd_559.packet_count,559);
      packet_count_check(port_count[560],env.pf_vf_mux_scbd_560.packet_count,560);
      packet_count_check(port_count[561],env.pf_vf_mux_scbd_561.packet_count,561);
      packet_count_check(port_count[562],env.pf_vf_mux_scbd_562.packet_count,562);
      packet_count_check(port_count[563],env.pf_vf_mux_scbd_563.packet_count,563);
      packet_count_check(port_count[564],env.pf_vf_mux_scbd_564.packet_count,564);
      packet_count_check(port_count[565],env.pf_vf_mux_scbd_565.packet_count,565);
      packet_count_check(port_count[566],env.pf_vf_mux_scbd_566.packet_count,566);
      packet_count_check(port_count[567],env.pf_vf_mux_scbd_567.packet_count,567);
      packet_count_check(port_count[568],env.pf_vf_mux_scbd_568.packet_count,568);
      packet_count_check(port_count[569],env.pf_vf_mux_scbd_569.packet_count,569);
      packet_count_check(port_count[570],env.pf_vf_mux_scbd_570.packet_count,570);
      packet_count_check(port_count[571],env.pf_vf_mux_scbd_571.packet_count,571);
      packet_count_check(port_count[572],env.pf_vf_mux_scbd_572.packet_count,572);
      packet_count_check(port_count[573],env.pf_vf_mux_scbd_573.packet_count,573);
      packet_count_check(port_count[574],env.pf_vf_mux_scbd_574.packet_count,574);
      packet_count_check(port_count[575],env.pf_vf_mux_scbd_575.packet_count,575);
      packet_count_check(port_count[576],env.pf_vf_mux_scbd_576.packet_count,576);
      packet_count_check(port_count[577],env.pf_vf_mux_scbd_577.packet_count,577);
      packet_count_check(port_count[578],env.pf_vf_mux_scbd_578.packet_count,578);
      packet_count_check(port_count[579],env.pf_vf_mux_scbd_579.packet_count,579);
      packet_count_check(port_count[580],env.pf_vf_mux_scbd_580.packet_count,580);
      packet_count_check(port_count[581],env.pf_vf_mux_scbd_581.packet_count,581);
      packet_count_check(port_count[582],env.pf_vf_mux_scbd_582.packet_count,582);
      packet_count_check(port_count[583],env.pf_vf_mux_scbd_583.packet_count,583);
      packet_count_check(port_count[584],env.pf_vf_mux_scbd_584.packet_count,584);
      packet_count_check(port_count[585],env.pf_vf_mux_scbd_585.packet_count,585);
      packet_count_check(port_count[586],env.pf_vf_mux_scbd_586.packet_count,586);
      packet_count_check(port_count[587],env.pf_vf_mux_scbd_587.packet_count,587);
      packet_count_check(port_count[588],env.pf_vf_mux_scbd_588.packet_count,588);
      packet_count_check(port_count[589],env.pf_vf_mux_scbd_589.packet_count,589);
      packet_count_check(port_count[590],env.pf_vf_mux_scbd_590.packet_count,590);
      packet_count_check(port_count[591],env.pf_vf_mux_scbd_591.packet_count,591);
      packet_count_check(port_count[592],env.pf_vf_mux_scbd_592.packet_count,592);
      packet_count_check(port_count[593],env.pf_vf_mux_scbd_593.packet_count,593);
      packet_count_check(port_count[594],env.pf_vf_mux_scbd_594.packet_count,594);
      packet_count_check(port_count[595],env.pf_vf_mux_scbd_595.packet_count,595);
      packet_count_check(port_count[596],env.pf_vf_mux_scbd_596.packet_count,596);
      packet_count_check(port_count[597],env.pf_vf_mux_scbd_597.packet_count,597);
      packet_count_check(port_count[598],env.pf_vf_mux_scbd_598.packet_count,598);
      packet_count_check(port_count[599],env.pf_vf_mux_scbd_599.packet_count,599);
      packet_count_check(port_count[600],env.pf_vf_mux_scbd_600.packet_count,600);
      packet_count_check(port_count[601],env.pf_vf_mux_scbd_601.packet_count,601);
      packet_count_check(port_count[602],env.pf_vf_mux_scbd_602.packet_count,602);
      packet_count_check(port_count[603],env.pf_vf_mux_scbd_603.packet_count,603);
      packet_count_check(port_count[604],env.pf_vf_mux_scbd_604.packet_count,604);
      packet_count_check(port_count[605],env.pf_vf_mux_scbd_605.packet_count,605);
      packet_count_check(port_count[606],env.pf_vf_mux_scbd_606.packet_count,606);
      packet_count_check(port_count[607],env.pf_vf_mux_scbd_607.packet_count,607);
      packet_count_check(port_count[608],env.pf_vf_mux_scbd_608.packet_count,608);
      packet_count_check(port_count[609],env.pf_vf_mux_scbd_609.packet_count,609);
      packet_count_check(port_count[610],env.pf_vf_mux_scbd_610.packet_count,610);
      packet_count_check(port_count[611],env.pf_vf_mux_scbd_611.packet_count,611);
      packet_count_check(port_count[612],env.pf_vf_mux_scbd_612.packet_count,612);
      packet_count_check(port_count[613],env.pf_vf_mux_scbd_613.packet_count,613);
      packet_count_check(port_count[614],env.pf_vf_mux_scbd_614.packet_count,614);
      packet_count_check(port_count[615],env.pf_vf_mux_scbd_615.packet_count,615);
      packet_count_check(port_count[616],env.pf_vf_mux_scbd_616.packet_count,616);
      packet_count_check(port_count[617],env.pf_vf_mux_scbd_617.packet_count,617);
      packet_count_check(port_count[618],env.pf_vf_mux_scbd_618.packet_count,618);
      packet_count_check(port_count[619],env.pf_vf_mux_scbd_619.packet_count,619);
      packet_count_check(port_count[620],env.pf_vf_mux_scbd_620.packet_count,620);
      packet_count_check(port_count[621],env.pf_vf_mux_scbd_621.packet_count,621);
      packet_count_check(port_count[622],env.pf_vf_mux_scbd_622.packet_count,622);
      packet_count_check(port_count[623],env.pf_vf_mux_scbd_623.packet_count,623);
      packet_count_check(port_count[624],env.pf_vf_mux_scbd_624.packet_count,624);
      packet_count_check(port_count[625],env.pf_vf_mux_scbd_625.packet_count,625);
      packet_count_check(port_count[626],env.pf_vf_mux_scbd_626.packet_count,626);
      packet_count_check(port_count[627],env.pf_vf_mux_scbd_627.packet_count,627);
      packet_count_check(port_count[628],env.pf_vf_mux_scbd_628.packet_count,628);
      packet_count_check(port_count[629],env.pf_vf_mux_scbd_629.packet_count,629);
      packet_count_check(port_count[630],env.pf_vf_mux_scbd_630.packet_count,630);
      packet_count_check(port_count[631],env.pf_vf_mux_scbd_631.packet_count,631);
      packet_count_check(port_count[632],env.pf_vf_mux_scbd_632.packet_count,632);
      packet_count_check(port_count[633],env.pf_vf_mux_scbd_633.packet_count,633);
      packet_count_check(port_count[634],env.pf_vf_mux_scbd_634.packet_count,634);
      packet_count_check(port_count[635],env.pf_vf_mux_scbd_635.packet_count,635);
      packet_count_check(port_count[636],env.pf_vf_mux_scbd_636.packet_count,636);
      packet_count_check(port_count[637],env.pf_vf_mux_scbd_637.packet_count,637);
      packet_count_check(port_count[638],env.pf_vf_mux_scbd_638.packet_count,638);
      packet_count_check(port_count[639],env.pf_vf_mux_scbd_639.packet_count,639);
      packet_count_check(port_count[640],env.pf_vf_mux_scbd_640.packet_count,640);
      packet_count_check(port_count[641],env.pf_vf_mux_scbd_641.packet_count,641);
      packet_count_check(port_count[642],env.pf_vf_mux_scbd_642.packet_count,642);
      packet_count_check(port_count[643],env.pf_vf_mux_scbd_643.packet_count,643);
      packet_count_check(port_count[644],env.pf_vf_mux_scbd_644.packet_count,644);
      packet_count_check(port_count[645],env.pf_vf_mux_scbd_645.packet_count,645);
      packet_count_check(port_count[646],env.pf_vf_mux_scbd_646.packet_count,646);
      packet_count_check(port_count[647],env.pf_vf_mux_scbd_647.packet_count,647);
      packet_count_check(port_count[648],env.pf_vf_mux_scbd_648.packet_count,648);
      packet_count_check(port_count[649],env.pf_vf_mux_scbd_649.packet_count,649);
      packet_count_check(port_count[650],env.pf_vf_mux_scbd_650.packet_count,650);
      packet_count_check(port_count[651],env.pf_vf_mux_scbd_651.packet_count,651);
      packet_count_check(port_count[652],env.pf_vf_mux_scbd_652.packet_count,652);
      packet_count_check(port_count[653],env.pf_vf_mux_scbd_653.packet_count,653);
      packet_count_check(port_count[654],env.pf_vf_mux_scbd_654.packet_count,654);
      packet_count_check(port_count[655],env.pf_vf_mux_scbd_655.packet_count,655);
      packet_count_check(port_count[656],env.pf_vf_mux_scbd_656.packet_count,656);
      packet_count_check(port_count[657],env.pf_vf_mux_scbd_657.packet_count,657);
      packet_count_check(port_count[658],env.pf_vf_mux_scbd_658.packet_count,658);
      packet_count_check(port_count[659],env.pf_vf_mux_scbd_659.packet_count,659);
      packet_count_check(port_count[660],env.pf_vf_mux_scbd_660.packet_count,660);
      packet_count_check(port_count[661],env.pf_vf_mux_scbd_661.packet_count,661);
      packet_count_check(port_count[662],env.pf_vf_mux_scbd_662.packet_count,662);
      packet_count_check(port_count[663],env.pf_vf_mux_scbd_663.packet_count,663);
      packet_count_check(port_count[664],env.pf_vf_mux_scbd_664.packet_count,664);
      packet_count_check(port_count[665],env.pf_vf_mux_scbd_665.packet_count,665);
      packet_count_check(port_count[666],env.pf_vf_mux_scbd_666.packet_count,666);
      packet_count_check(port_count[667],env.pf_vf_mux_scbd_667.packet_count,667);
      packet_count_check(port_count[668],env.pf_vf_mux_scbd_668.packet_count,668);
      packet_count_check(port_count[669],env.pf_vf_mux_scbd_669.packet_count,669);
      packet_count_check(port_count[670],env.pf_vf_mux_scbd_670.packet_count,670);
      packet_count_check(port_count[671],env.pf_vf_mux_scbd_671.packet_count,671);
      packet_count_check(port_count[672],env.pf_vf_mux_scbd_672.packet_count,672);
      packet_count_check(port_count[673],env.pf_vf_mux_scbd_673.packet_count,673);
      packet_count_check(port_count[674],env.pf_vf_mux_scbd_674.packet_count,674);
      packet_count_check(port_count[675],env.pf_vf_mux_scbd_675.packet_count,675);
      packet_count_check(port_count[676],env.pf_vf_mux_scbd_676.packet_count,676);
      packet_count_check(port_count[677],env.pf_vf_mux_scbd_677.packet_count,677);
      packet_count_check(port_count[678],env.pf_vf_mux_scbd_678.packet_count,678);
      packet_count_check(port_count[679],env.pf_vf_mux_scbd_679.packet_count,679);
      packet_count_check(port_count[680],env.pf_vf_mux_scbd_680.packet_count,680);
      packet_count_check(port_count[681],env.pf_vf_mux_scbd_681.packet_count,681);
      packet_count_check(port_count[682],env.pf_vf_mux_scbd_682.packet_count,682);
      packet_count_check(port_count[683],env.pf_vf_mux_scbd_683.packet_count,683);
      packet_count_check(port_count[684],env.pf_vf_mux_scbd_684.packet_count,684);
      packet_count_check(port_count[685],env.pf_vf_mux_scbd_685.packet_count,685);
      packet_count_check(port_count[686],env.pf_vf_mux_scbd_686.packet_count,686);
      packet_count_check(port_count[687],env.pf_vf_mux_scbd_687.packet_count,687);
      packet_count_check(port_count[688],env.pf_vf_mux_scbd_688.packet_count,688);
      packet_count_check(port_count[689],env.pf_vf_mux_scbd_689.packet_count,689);
      packet_count_check(port_count[690],env.pf_vf_mux_scbd_690.packet_count,690);
      packet_count_check(port_count[691],env.pf_vf_mux_scbd_691.packet_count,691);
      packet_count_check(port_count[692],env.pf_vf_mux_scbd_692.packet_count,692);
      packet_count_check(port_count[693],env.pf_vf_mux_scbd_693.packet_count,693);
      packet_count_check(port_count[694],env.pf_vf_mux_scbd_694.packet_count,694);
      packet_count_check(port_count[695],env.pf_vf_mux_scbd_695.packet_count,695);
      packet_count_check(port_count[696],env.pf_vf_mux_scbd_696.packet_count,696);
      packet_count_check(port_count[697],env.pf_vf_mux_scbd_697.packet_count,697);
      packet_count_check(port_count[698],env.pf_vf_mux_scbd_698.packet_count,698);
      packet_count_check(port_count[699],env.pf_vf_mux_scbd_699.packet_count,699);
      packet_count_check(port_count[700],env.pf_vf_mux_scbd_700.packet_count,700);
      packet_count_check(port_count[701],env.pf_vf_mux_scbd_701.packet_count,701);
      packet_count_check(port_count[702],env.pf_vf_mux_scbd_702.packet_count,702);
      packet_count_check(port_count[703],env.pf_vf_mux_scbd_703.packet_count,703);
      packet_count_check(port_count[704],env.pf_vf_mux_scbd_704.packet_count,704);
      packet_count_check(port_count[705],env.pf_vf_mux_scbd_705.packet_count,705);
      packet_count_check(port_count[706],env.pf_vf_mux_scbd_706.packet_count,706);
      packet_count_check(port_count[707],env.pf_vf_mux_scbd_707.packet_count,707);
      packet_count_check(port_count[708],env.pf_vf_mux_scbd_708.packet_count,708);
      packet_count_check(port_count[709],env.pf_vf_mux_scbd_709.packet_count,709);
      packet_count_check(port_count[710],env.pf_vf_mux_scbd_710.packet_count,710);
      packet_count_check(port_count[711],env.pf_vf_mux_scbd_711.packet_count,711);
      packet_count_check(port_count[712],env.pf_vf_mux_scbd_712.packet_count,712);
      packet_count_check(port_count[713],env.pf_vf_mux_scbd_713.packet_count,713);
      packet_count_check(port_count[714],env.pf_vf_mux_scbd_714.packet_count,714);
      packet_count_check(port_count[715],env.pf_vf_mux_scbd_715.packet_count,715);
      packet_count_check(port_count[716],env.pf_vf_mux_scbd_716.packet_count,716);
      packet_count_check(port_count[717],env.pf_vf_mux_scbd_717.packet_count,717);
      packet_count_check(port_count[718],env.pf_vf_mux_scbd_718.packet_count,718);
      packet_count_check(port_count[719],env.pf_vf_mux_scbd_719.packet_count,719);
      packet_count_check(port_count[720],env.pf_vf_mux_scbd_720.packet_count,720);
      packet_count_check(port_count[721],env.pf_vf_mux_scbd_721.packet_count,721);
      packet_count_check(port_count[722],env.pf_vf_mux_scbd_722.packet_count,722);
      packet_count_check(port_count[723],env.pf_vf_mux_scbd_723.packet_count,723);
      packet_count_check(port_count[724],env.pf_vf_mux_scbd_724.packet_count,724);
      packet_count_check(port_count[725],env.pf_vf_mux_scbd_725.packet_count,725);
      packet_count_check(port_count[726],env.pf_vf_mux_scbd_726.packet_count,726);
      packet_count_check(port_count[727],env.pf_vf_mux_scbd_727.packet_count,727);
      packet_count_check(port_count[728],env.pf_vf_mux_scbd_728.packet_count,728);
      packet_count_check(port_count[729],env.pf_vf_mux_scbd_729.packet_count,729);
      packet_count_check(port_count[730],env.pf_vf_mux_scbd_730.packet_count,730);
      packet_count_check(port_count[731],env.pf_vf_mux_scbd_731.packet_count,731);
      packet_count_check(port_count[732],env.pf_vf_mux_scbd_732.packet_count,732);
      packet_count_check(port_count[733],env.pf_vf_mux_scbd_733.packet_count,733);
      packet_count_check(port_count[734],env.pf_vf_mux_scbd_734.packet_count,734);
      packet_count_check(port_count[735],env.pf_vf_mux_scbd_735.packet_count,735);
      packet_count_check(port_count[736],env.pf_vf_mux_scbd_736.packet_count,736);
      packet_count_check(port_count[737],env.pf_vf_mux_scbd_737.packet_count,737);
      packet_count_check(port_count[738],env.pf_vf_mux_scbd_738.packet_count,738);
      packet_count_check(port_count[739],env.pf_vf_mux_scbd_739.packet_count,739);
      packet_count_check(port_count[740],env.pf_vf_mux_scbd_740.packet_count,740);
      packet_count_check(port_count[741],env.pf_vf_mux_scbd_741.packet_count,741);
      packet_count_check(port_count[742],env.pf_vf_mux_scbd_742.packet_count,742);
      packet_count_check(port_count[743],env.pf_vf_mux_scbd_743.packet_count,743);
      packet_count_check(port_count[744],env.pf_vf_mux_scbd_744.packet_count,744);
      packet_count_check(port_count[745],env.pf_vf_mux_scbd_745.packet_count,745);
      packet_count_check(port_count[746],env.pf_vf_mux_scbd_746.packet_count,746);
      packet_count_check(port_count[747],env.pf_vf_mux_scbd_747.packet_count,747);
      packet_count_check(port_count[748],env.pf_vf_mux_scbd_748.packet_count,748);
      packet_count_check(port_count[749],env.pf_vf_mux_scbd_749.packet_count,749);
      packet_count_check(port_count[750],env.pf_vf_mux_scbd_750.packet_count,750);
      packet_count_check(port_count[751],env.pf_vf_mux_scbd_751.packet_count,751);
      packet_count_check(port_count[752],env.pf_vf_mux_scbd_752.packet_count,752);
      packet_count_check(port_count[753],env.pf_vf_mux_scbd_753.packet_count,753);
      packet_count_check(port_count[754],env.pf_vf_mux_scbd_754.packet_count,754);
      packet_count_check(port_count[755],env.pf_vf_mux_scbd_755.packet_count,755);
      packet_count_check(port_count[756],env.pf_vf_mux_scbd_756.packet_count,756);
      packet_count_check(port_count[757],env.pf_vf_mux_scbd_757.packet_count,757);
      packet_count_check(port_count[758],env.pf_vf_mux_scbd_758.packet_count,758);
      packet_count_check(port_count[759],env.pf_vf_mux_scbd_759.packet_count,759);
      packet_count_check(port_count[760],env.pf_vf_mux_scbd_760.packet_count,760);
      packet_count_check(port_count[761],env.pf_vf_mux_scbd_761.packet_count,761);
      packet_count_check(port_count[762],env.pf_vf_mux_scbd_762.packet_count,762);
      packet_count_check(port_count[763],env.pf_vf_mux_scbd_763.packet_count,763);
      packet_count_check(port_count[764],env.pf_vf_mux_scbd_764.packet_count,764);
      packet_count_check(port_count[765],env.pf_vf_mux_scbd_765.packet_count,765);
      packet_count_check(port_count[766],env.pf_vf_mux_scbd_766.packet_count,766);
      packet_count_check(port_count[767],env.pf_vf_mux_scbd_767.packet_count,767);
      packet_count_check(port_count[768],env.pf_vf_mux_scbd_768.packet_count,768);
      packet_count_check(port_count[769],env.pf_vf_mux_scbd_769.packet_count,769);
      packet_count_check(port_count[770],env.pf_vf_mux_scbd_770.packet_count,770);
      packet_count_check(port_count[771],env.pf_vf_mux_scbd_771.packet_count,771);
      packet_count_check(port_count[772],env.pf_vf_mux_scbd_772.packet_count,772);
      packet_count_check(port_count[773],env.pf_vf_mux_scbd_773.packet_count,773);
      packet_count_check(port_count[774],env.pf_vf_mux_scbd_774.packet_count,774);
      packet_count_check(port_count[775],env.pf_vf_mux_scbd_775.packet_count,775);
      packet_count_check(port_count[776],env.pf_vf_mux_scbd_776.packet_count,776);
      packet_count_check(port_count[777],env.pf_vf_mux_scbd_777.packet_count,777);
      packet_count_check(port_count[778],env.pf_vf_mux_scbd_778.packet_count,778);
      packet_count_check(port_count[779],env.pf_vf_mux_scbd_779.packet_count,779);
      packet_count_check(port_count[780],env.pf_vf_mux_scbd_780.packet_count,780);
      packet_count_check(port_count[781],env.pf_vf_mux_scbd_781.packet_count,781);
      packet_count_check(port_count[782],env.pf_vf_mux_scbd_782.packet_count,782);
      packet_count_check(port_count[783],env.pf_vf_mux_scbd_783.packet_count,783);
      packet_count_check(port_count[784],env.pf_vf_mux_scbd_784.packet_count,784);
      packet_count_check(port_count[785],env.pf_vf_mux_scbd_785.packet_count,785);
      packet_count_check(port_count[786],env.pf_vf_mux_scbd_786.packet_count,786);
      packet_count_check(port_count[787],env.pf_vf_mux_scbd_787.packet_count,787);
      packet_count_check(port_count[788],env.pf_vf_mux_scbd_788.packet_count,788);
      packet_count_check(port_count[789],env.pf_vf_mux_scbd_789.packet_count,789);
      packet_count_check(port_count[790],env.pf_vf_mux_scbd_790.packet_count,790);
      packet_count_check(port_count[791],env.pf_vf_mux_scbd_791.packet_count,791);
      packet_count_check(port_count[792],env.pf_vf_mux_scbd_792.packet_count,792);
      packet_count_check(port_count[793],env.pf_vf_mux_scbd_793.packet_count,793);
      packet_count_check(port_count[794],env.pf_vf_mux_scbd_794.packet_count,794);
      packet_count_check(port_count[795],env.pf_vf_mux_scbd_795.packet_count,795);
      packet_count_check(port_count[796],env.pf_vf_mux_scbd_796.packet_count,796);
      packet_count_check(port_count[797],env.pf_vf_mux_scbd_797.packet_count,797);
      packet_count_check(port_count[798],env.pf_vf_mux_scbd_798.packet_count,798);
      packet_count_check(port_count[799],env.pf_vf_mux_scbd_799.packet_count,799);
      packet_count_check(port_count[800],env.pf_vf_mux_scbd_800.packet_count,800);
      packet_count_check(port_count[801],env.pf_vf_mux_scbd_801.packet_count,801);
      packet_count_check(port_count[802],env.pf_vf_mux_scbd_802.packet_count,802);
      packet_count_check(port_count[803],env.pf_vf_mux_scbd_803.packet_count,803);
      packet_count_check(port_count[804],env.pf_vf_mux_scbd_804.packet_count,804);
      packet_count_check(port_count[805],env.pf_vf_mux_scbd_805.packet_count,805);
      packet_count_check(port_count[806],env.pf_vf_mux_scbd_806.packet_count,806);
      packet_count_check(port_count[807],env.pf_vf_mux_scbd_807.packet_count,807);
      packet_count_check(port_count[808],env.pf_vf_mux_scbd_808.packet_count,808);
      packet_count_check(port_count[809],env.pf_vf_mux_scbd_809.packet_count,809);
      packet_count_check(port_count[810],env.pf_vf_mux_scbd_810.packet_count,810);
      packet_count_check(port_count[811],env.pf_vf_mux_scbd_811.packet_count,811);
      packet_count_check(port_count[812],env.pf_vf_mux_scbd_812.packet_count,812);
      packet_count_check(port_count[813],env.pf_vf_mux_scbd_813.packet_count,813);
      packet_count_check(port_count[814],env.pf_vf_mux_scbd_814.packet_count,814);
      packet_count_check(port_count[815],env.pf_vf_mux_scbd_815.packet_count,815);
      packet_count_check(port_count[816],env.pf_vf_mux_scbd_816.packet_count,816);
      packet_count_check(port_count[817],env.pf_vf_mux_scbd_817.packet_count,817);
      packet_count_check(port_count[818],env.pf_vf_mux_scbd_818.packet_count,818);
      packet_count_check(port_count[819],env.pf_vf_mux_scbd_819.packet_count,819);
      packet_count_check(port_count[820],env.pf_vf_mux_scbd_820.packet_count,820);
      packet_count_check(port_count[821],env.pf_vf_mux_scbd_821.packet_count,821);
      packet_count_check(port_count[822],env.pf_vf_mux_scbd_822.packet_count,822);
      packet_count_check(port_count[823],env.pf_vf_mux_scbd_823.packet_count,823);
      packet_count_check(port_count[824],env.pf_vf_mux_scbd_824.packet_count,824);
      packet_count_check(port_count[825],env.pf_vf_mux_scbd_825.packet_count,825);
      packet_count_check(port_count[826],env.pf_vf_mux_scbd_826.packet_count,826);
      packet_count_check(port_count[827],env.pf_vf_mux_scbd_827.packet_count,827);
      packet_count_check(port_count[828],env.pf_vf_mux_scbd_828.packet_count,828);
      packet_count_check(port_count[829],env.pf_vf_mux_scbd_829.packet_count,829);
      packet_count_check(port_count[830],env.pf_vf_mux_scbd_830.packet_count,830);
      packet_count_check(port_count[831],env.pf_vf_mux_scbd_831.packet_count,831);
      packet_count_check(port_count[832],env.pf_vf_mux_scbd_832.packet_count,832);
      packet_count_check(port_count[833],env.pf_vf_mux_scbd_833.packet_count,833);
      packet_count_check(port_count[834],env.pf_vf_mux_scbd_834.packet_count,834);
      packet_count_check(port_count[835],env.pf_vf_mux_scbd_835.packet_count,835);
      packet_count_check(port_count[836],env.pf_vf_mux_scbd_836.packet_count,836);
      packet_count_check(port_count[837],env.pf_vf_mux_scbd_837.packet_count,837);
      packet_count_check(port_count[838],env.pf_vf_mux_scbd_838.packet_count,838);
      packet_count_check(port_count[839],env.pf_vf_mux_scbd_839.packet_count,839);
      packet_count_check(port_count[840],env.pf_vf_mux_scbd_840.packet_count,840);
      packet_count_check(port_count[841],env.pf_vf_mux_scbd_841.packet_count,841);
      packet_count_check(port_count[842],env.pf_vf_mux_scbd_842.packet_count,842);
      packet_count_check(port_count[843],env.pf_vf_mux_scbd_843.packet_count,843);
      packet_count_check(port_count[844],env.pf_vf_mux_scbd_844.packet_count,844);
      packet_count_check(port_count[845],env.pf_vf_mux_scbd_845.packet_count,845);
      packet_count_check(port_count[846],env.pf_vf_mux_scbd_846.packet_count,846);
      packet_count_check(port_count[847],env.pf_vf_mux_scbd_847.packet_count,847);
      packet_count_check(port_count[848],env.pf_vf_mux_scbd_848.packet_count,848);
      packet_count_check(port_count[849],env.pf_vf_mux_scbd_849.packet_count,849);
      packet_count_check(port_count[850],env.pf_vf_mux_scbd_850.packet_count,850);
      packet_count_check(port_count[851],env.pf_vf_mux_scbd_851.packet_count,851);
      packet_count_check(port_count[852],env.pf_vf_mux_scbd_852.packet_count,852);
      packet_count_check(port_count[853],env.pf_vf_mux_scbd_853.packet_count,853);
      packet_count_check(port_count[854],env.pf_vf_mux_scbd_854.packet_count,854);
      packet_count_check(port_count[855],env.pf_vf_mux_scbd_855.packet_count,855);
      packet_count_check(port_count[856],env.pf_vf_mux_scbd_856.packet_count,856);
      packet_count_check(port_count[857],env.pf_vf_mux_scbd_857.packet_count,857);
      packet_count_check(port_count[858],env.pf_vf_mux_scbd_858.packet_count,858);
      packet_count_check(port_count[859],env.pf_vf_mux_scbd_859.packet_count,859);
      packet_count_check(port_count[860],env.pf_vf_mux_scbd_860.packet_count,860);
      packet_count_check(port_count[861],env.pf_vf_mux_scbd_861.packet_count,861);
      packet_count_check(port_count[862],env.pf_vf_mux_scbd_862.packet_count,862);
      packet_count_check(port_count[863],env.pf_vf_mux_scbd_863.packet_count,863);
      packet_count_check(port_count[864],env.pf_vf_mux_scbd_864.packet_count,864);
      packet_count_check(port_count[865],env.pf_vf_mux_scbd_865.packet_count,865);
      packet_count_check(port_count[866],env.pf_vf_mux_scbd_866.packet_count,866);
      packet_count_check(port_count[867],env.pf_vf_mux_scbd_867.packet_count,867);
      packet_count_check(port_count[868],env.pf_vf_mux_scbd_868.packet_count,868);
      packet_count_check(port_count[869],env.pf_vf_mux_scbd_869.packet_count,869);
      packet_count_check(port_count[870],env.pf_vf_mux_scbd_870.packet_count,870);
      packet_count_check(port_count[871],env.pf_vf_mux_scbd_871.packet_count,871);
      packet_count_check(port_count[872],env.pf_vf_mux_scbd_872.packet_count,872);
      packet_count_check(port_count[873],env.pf_vf_mux_scbd_873.packet_count,873);
      packet_count_check(port_count[874],env.pf_vf_mux_scbd_874.packet_count,874);
      packet_count_check(port_count[875],env.pf_vf_mux_scbd_875.packet_count,875);
      packet_count_check(port_count[876],env.pf_vf_mux_scbd_876.packet_count,876);
      packet_count_check(port_count[877],env.pf_vf_mux_scbd_877.packet_count,877);
      packet_count_check(port_count[878],env.pf_vf_mux_scbd_878.packet_count,878);
      packet_count_check(port_count[879],env.pf_vf_mux_scbd_879.packet_count,879);
      packet_count_check(port_count[880],env.pf_vf_mux_scbd_880.packet_count,880);
      packet_count_check(port_count[881],env.pf_vf_mux_scbd_881.packet_count,881);
      packet_count_check(port_count[882],env.pf_vf_mux_scbd_882.packet_count,882);
      packet_count_check(port_count[883],env.pf_vf_mux_scbd_883.packet_count,883);
      packet_count_check(port_count[884],env.pf_vf_mux_scbd_884.packet_count,884);
      packet_count_check(port_count[885],env.pf_vf_mux_scbd_885.packet_count,885);
      packet_count_check(port_count[886],env.pf_vf_mux_scbd_886.packet_count,886);
      packet_count_check(port_count[887],env.pf_vf_mux_scbd_887.packet_count,887);
      packet_count_check(port_count[888],env.pf_vf_mux_scbd_888.packet_count,888);
      packet_count_check(port_count[889],env.pf_vf_mux_scbd_889.packet_count,889);
      packet_count_check(port_count[890],env.pf_vf_mux_scbd_890.packet_count,890);
      packet_count_check(port_count[891],env.pf_vf_mux_scbd_891.packet_count,891);
      packet_count_check(port_count[892],env.pf_vf_mux_scbd_892.packet_count,892);
      packet_count_check(port_count[893],env.pf_vf_mux_scbd_893.packet_count,893);
      packet_count_check(port_count[894],env.pf_vf_mux_scbd_894.packet_count,894);
      packet_count_check(port_count[895],env.pf_vf_mux_scbd_895.packet_count,895);
      packet_count_check(port_count[896],env.pf_vf_mux_scbd_896.packet_count,896);
      packet_count_check(port_count[897],env.pf_vf_mux_scbd_897.packet_count,897);
      packet_count_check(port_count[898],env.pf_vf_mux_scbd_898.packet_count,898);
      packet_count_check(port_count[899],env.pf_vf_mux_scbd_899.packet_count,899);
      packet_count_check(port_count[900],env.pf_vf_mux_scbd_900.packet_count,900);
      packet_count_check(port_count[901],env.pf_vf_mux_scbd_901.packet_count,901);
      packet_count_check(port_count[902],env.pf_vf_mux_scbd_902.packet_count,902);
      packet_count_check(port_count[903],env.pf_vf_mux_scbd_903.packet_count,903);
      packet_count_check(port_count[904],env.pf_vf_mux_scbd_904.packet_count,904);
      packet_count_check(port_count[905],env.pf_vf_mux_scbd_905.packet_count,905);
      packet_count_check(port_count[906],env.pf_vf_mux_scbd_906.packet_count,906);
      packet_count_check(port_count[907],env.pf_vf_mux_scbd_907.packet_count,907);
      packet_count_check(port_count[908],env.pf_vf_mux_scbd_908.packet_count,908);
      packet_count_check(port_count[909],env.pf_vf_mux_scbd_909.packet_count,909);
      packet_count_check(port_count[910],env.pf_vf_mux_scbd_910.packet_count,910);
      packet_count_check(port_count[911],env.pf_vf_mux_scbd_911.packet_count,911);
      packet_count_check(port_count[912],env.pf_vf_mux_scbd_912.packet_count,912);
      packet_count_check(port_count[913],env.pf_vf_mux_scbd_913.packet_count,913);
      packet_count_check(port_count[914],env.pf_vf_mux_scbd_914.packet_count,914);
      packet_count_check(port_count[915],env.pf_vf_mux_scbd_915.packet_count,915);
      packet_count_check(port_count[916],env.pf_vf_mux_scbd_916.packet_count,916);
      packet_count_check(port_count[917],env.pf_vf_mux_scbd_917.packet_count,917);
      packet_count_check(port_count[918],env.pf_vf_mux_scbd_918.packet_count,918);
      packet_count_check(port_count[919],env.pf_vf_mux_scbd_919.packet_count,919);
      packet_count_check(port_count[920],env.pf_vf_mux_scbd_920.packet_count,920);
      packet_count_check(port_count[921],env.pf_vf_mux_scbd_921.packet_count,921);
      packet_count_check(port_count[922],env.pf_vf_mux_scbd_922.packet_count,922);
      packet_count_check(port_count[923],env.pf_vf_mux_scbd_923.packet_count,923);
      packet_count_check(port_count[924],env.pf_vf_mux_scbd_924.packet_count,924);
      packet_count_check(port_count[925],env.pf_vf_mux_scbd_925.packet_count,925);
      packet_count_check(port_count[926],env.pf_vf_mux_scbd_926.packet_count,926);
      packet_count_check(port_count[927],env.pf_vf_mux_scbd_927.packet_count,927);
      packet_count_check(port_count[928],env.pf_vf_mux_scbd_928.packet_count,928);
      packet_count_check(port_count[929],env.pf_vf_mux_scbd_929.packet_count,929);
      packet_count_check(port_count[930],env.pf_vf_mux_scbd_930.packet_count,930);
      packet_count_check(port_count[931],env.pf_vf_mux_scbd_931.packet_count,931);
      packet_count_check(port_count[932],env.pf_vf_mux_scbd_932.packet_count,932);
      packet_count_check(port_count[933],env.pf_vf_mux_scbd_933.packet_count,933);
      packet_count_check(port_count[934],env.pf_vf_mux_scbd_934.packet_count,934);
      packet_count_check(port_count[935],env.pf_vf_mux_scbd_935.packet_count,935);
      packet_count_check(port_count[936],env.pf_vf_mux_scbd_936.packet_count,936);
      packet_count_check(port_count[937],env.pf_vf_mux_scbd_937.packet_count,937);
      packet_count_check(port_count[938],env.pf_vf_mux_scbd_938.packet_count,938);
      packet_count_check(port_count[939],env.pf_vf_mux_scbd_939.packet_count,939);
      packet_count_check(port_count[940],env.pf_vf_mux_scbd_940.packet_count,940);
      packet_count_check(port_count[941],env.pf_vf_mux_scbd_941.packet_count,941);
      packet_count_check(port_count[942],env.pf_vf_mux_scbd_942.packet_count,942);
      packet_count_check(port_count[943],env.pf_vf_mux_scbd_943.packet_count,943);
      packet_count_check(port_count[944],env.pf_vf_mux_scbd_944.packet_count,944);
      packet_count_check(port_count[945],env.pf_vf_mux_scbd_945.packet_count,945);
      packet_count_check(port_count[946],env.pf_vf_mux_scbd_946.packet_count,946);
      packet_count_check(port_count[947],env.pf_vf_mux_scbd_947.packet_count,947);
      packet_count_check(port_count[948],env.pf_vf_mux_scbd_948.packet_count,948);
      packet_count_check(port_count[949],env.pf_vf_mux_scbd_949.packet_count,949);
      packet_count_check(port_count[950],env.pf_vf_mux_scbd_950.packet_count,950);
      packet_count_check(port_count[951],env.pf_vf_mux_scbd_951.packet_count,951);
      packet_count_check(port_count[952],env.pf_vf_mux_scbd_952.packet_count,952);
      packet_count_check(port_count[953],env.pf_vf_mux_scbd_953.packet_count,953);
      packet_count_check(port_count[954],env.pf_vf_mux_scbd_954.packet_count,954);
      packet_count_check(port_count[955],env.pf_vf_mux_scbd_955.packet_count,955);
      packet_count_check(port_count[956],env.pf_vf_mux_scbd_956.packet_count,956);
      packet_count_check(port_count[957],env.pf_vf_mux_scbd_957.packet_count,957);
      packet_count_check(port_count[958],env.pf_vf_mux_scbd_958.packet_count,958);
      packet_count_check(port_count[959],env.pf_vf_mux_scbd_959.packet_count,959);
      packet_count_check(port_count[960],env.pf_vf_mux_scbd_960.packet_count,960);
      packet_count_check(port_count[961],env.pf_vf_mux_scbd_961.packet_count,961);
      packet_count_check(port_count[962],env.pf_vf_mux_scbd_962.packet_count,962);
      packet_count_check(port_count[963],env.pf_vf_mux_scbd_963.packet_count,963);
      packet_count_check(port_count[964],env.pf_vf_mux_scbd_964.packet_count,964);
      packet_count_check(port_count[965],env.pf_vf_mux_scbd_965.packet_count,965);
      packet_count_check(port_count[966],env.pf_vf_mux_scbd_966.packet_count,966);
      packet_count_check(port_count[967],env.pf_vf_mux_scbd_967.packet_count,967);
      packet_count_check(port_count[968],env.pf_vf_mux_scbd_968.packet_count,968);
      packet_count_check(port_count[969],env.pf_vf_mux_scbd_969.packet_count,969);
      packet_count_check(port_count[970],env.pf_vf_mux_scbd_970.packet_count,970);
      packet_count_check(port_count[971],env.pf_vf_mux_scbd_971.packet_count,971);
      packet_count_check(port_count[972],env.pf_vf_mux_scbd_972.packet_count,972);
      packet_count_check(port_count[973],env.pf_vf_mux_scbd_973.packet_count,973);
      packet_count_check(port_count[974],env.pf_vf_mux_scbd_974.packet_count,974);
      packet_count_check(port_count[975],env.pf_vf_mux_scbd_975.packet_count,975);
      packet_count_check(port_count[976],env.pf_vf_mux_scbd_976.packet_count,976);
      packet_count_check(port_count[977],env.pf_vf_mux_scbd_977.packet_count,977);
      packet_count_check(port_count[978],env.pf_vf_mux_scbd_978.packet_count,978);
      packet_count_check(port_count[979],env.pf_vf_mux_scbd_979.packet_count,979);
      packet_count_check(port_count[980],env.pf_vf_mux_scbd_980.packet_count,980);
      packet_count_check(port_count[981],env.pf_vf_mux_scbd_981.packet_count,981);
      packet_count_check(port_count[982],env.pf_vf_mux_scbd_982.packet_count,982);
      packet_count_check(port_count[983],env.pf_vf_mux_scbd_983.packet_count,983);
      packet_count_check(port_count[984],env.pf_vf_mux_scbd_984.packet_count,984);
      packet_count_check(port_count[985],env.pf_vf_mux_scbd_985.packet_count,985);
      packet_count_check(port_count[986],env.pf_vf_mux_scbd_986.packet_count,986);
      packet_count_check(port_count[987],env.pf_vf_mux_scbd_987.packet_count,987);
      packet_count_check(port_count[988],env.pf_vf_mux_scbd_988.packet_count,988);
      packet_count_check(port_count[989],env.pf_vf_mux_scbd_989.packet_count,989);
      packet_count_check(port_count[990],env.pf_vf_mux_scbd_990.packet_count,990);
      packet_count_check(port_count[991],env.pf_vf_mux_scbd_991.packet_count,991);
      packet_count_check(port_count[992],env.pf_vf_mux_scbd_992.packet_count,992);
      packet_count_check(port_count[993],env.pf_vf_mux_scbd_993.packet_count,993);
      packet_count_check(port_count[994],env.pf_vf_mux_scbd_994.packet_count,994);
      packet_count_check(port_count[995],env.pf_vf_mux_scbd_995.packet_count,995);
      packet_count_check(port_count[996],env.pf_vf_mux_scbd_996.packet_count,996);
      packet_count_check(port_count[997],env.pf_vf_mux_scbd_997.packet_count,997);
      packet_count_check(port_count[998],env.pf_vf_mux_scbd_998.packet_count,998);
      packet_count_check(port_count[999],env.pf_vf_mux_scbd_999.packet_count,999);
      packet_count_check(port_count[1000],env.pf_vf_mux_scbd_1000.packet_count,1000);
      packet_count_check(port_count[1001],env.pf_vf_mux_scbd_1001.packet_count,1001);
      packet_count_check(port_count[1002],env.pf_vf_mux_scbd_1002.packet_count,1002);
      packet_count_check(port_count[1003],env.pf_vf_mux_scbd_1003.packet_count,1003);
      packet_count_check(port_count[1004],env.pf_vf_mux_scbd_1004.packet_count,1004);
      packet_count_check(port_count[1005],env.pf_vf_mux_scbd_1005.packet_count,1005);
      packet_count_check(port_count[1006],env.pf_vf_mux_scbd_1006.packet_count,1006);
      packet_count_check(port_count[1007],env.pf_vf_mux_scbd_1007.packet_count,1007);
      packet_count_check(port_count[1008],env.pf_vf_mux_scbd_1008.packet_count,1008);
      packet_count_check(port_count[1009],env.pf_vf_mux_scbd_1009.packet_count,1009);
      packet_count_check(port_count[1010],env.pf_vf_mux_scbd_1010.packet_count,1010);
      packet_count_check(port_count[1011],env.pf_vf_mux_scbd_1011.packet_count,1011);
      packet_count_check(port_count[1012],env.pf_vf_mux_scbd_1012.packet_count,1012);
      packet_count_check(port_count[1013],env.pf_vf_mux_scbd_1013.packet_count,1013);
      packet_count_check(port_count[1014],env.pf_vf_mux_scbd_1014.packet_count,1014);
      packet_count_check(port_count[1015],env.pf_vf_mux_scbd_1015.packet_count,1015);
      packet_count_check(port_count[1016],env.pf_vf_mux_scbd_1016.packet_count,1016);
      packet_count_check(port_count[1017],env.pf_vf_mux_scbd_1017.packet_count,1017);
      packet_count_check(port_count[1018],env.pf_vf_mux_scbd_1018.packet_count,1018);
      packet_count_check(port_count[1019],env.pf_vf_mux_scbd_1019.packet_count,1019);
      packet_count_check(port_count[1020],env.pf_vf_mux_scbd_1020.packet_count,1020);
      packet_count_check(port_count[1021],env.pf_vf_mux_scbd_1021.packet_count,1021);
      packet_count_check(port_count[1022],env.pf_vf_mux_scbd_1022.packet_count,1022);
      packet_count_check(port_count[1023],env.pf_vf_mux_scbd_1023.packet_count,1023);
      packet_count_check(port_count[1024],env.pf_vf_mux_scbd_1024.packet_count,1024);
      packet_count_check(port_count[1025],env.pf_vf_mux_scbd_1025.packet_count,1025);
      packet_count_check(port_count[1026],env.pf_vf_mux_scbd_1026.packet_count,1026);
      packet_count_check(port_count[1027],env.pf_vf_mux_scbd_1027.packet_count,1027);
      packet_count_check(port_count[1028],env.pf_vf_mux_scbd_1028.packet_count,1028);
      packet_count_check(port_count[1029],env.pf_vf_mux_scbd_1029.packet_count,1029);
      packet_count_check(port_count[1030],env.pf_vf_mux_scbd_1030.packet_count,1030);
      packet_count_check(port_count[1031],env.pf_vf_mux_scbd_1031.packet_count,1031);
      packet_count_check(port_count[1032],env.pf_vf_mux_scbd_1032.packet_count,1032);
      packet_count_check(port_count[1033],env.pf_vf_mux_scbd_1033.packet_count,1033);
      packet_count_check(port_count[1034],env.pf_vf_mux_scbd_1034.packet_count,1034);
      packet_count_check(port_count[1035],env.pf_vf_mux_scbd_1035.packet_count,1035);
      packet_count_check(port_count[1036],env.pf_vf_mux_scbd_1036.packet_count,1036);
      packet_count_check(port_count[1037],env.pf_vf_mux_scbd_1037.packet_count,1037);
      packet_count_check(port_count[1038],env.pf_vf_mux_scbd_1038.packet_count,1038);
      packet_count_check(port_count[1039],env.pf_vf_mux_scbd_1039.packet_count,1039);
      packet_count_check(port_count[1040],env.pf_vf_mux_scbd_1040.packet_count,1040);
      packet_count_check(port_count[1041],env.pf_vf_mux_scbd_1041.packet_count,1041);
      packet_count_check(port_count[1042],env.pf_vf_mux_scbd_1042.packet_count,1042);
      packet_count_check(port_count[1043],env.pf_vf_mux_scbd_1043.packet_count,1043);
      packet_count_check(port_count[1044],env.pf_vf_mux_scbd_1044.packet_count,1044);
      packet_count_check(port_count[1045],env.pf_vf_mux_scbd_1045.packet_count,1045);
      packet_count_check(port_count[1046],env.pf_vf_mux_scbd_1046.packet_count,1046);
      packet_count_check(port_count[1047],env.pf_vf_mux_scbd_1047.packet_count,1047);
      packet_count_check(port_count[1048],env.pf_vf_mux_scbd_1048.packet_count,1048);
      packet_count_check(port_count[1049],env.pf_vf_mux_scbd_1049.packet_count,1049);
      packet_count_check(port_count[1050],env.pf_vf_mux_scbd_1050.packet_count,1050);
      packet_count_check(port_count[1051],env.pf_vf_mux_scbd_1051.packet_count,1051);
      packet_count_check(port_count[1052],env.pf_vf_mux_scbd_1052.packet_count,1052);
      packet_count_check(port_count[1053],env.pf_vf_mux_scbd_1053.packet_count,1053);
      packet_count_check(port_count[1054],env.pf_vf_mux_scbd_1054.packet_count,1054);
      packet_count_check(port_count[1055],env.pf_vf_mux_scbd_1055.packet_count,1055);
      packet_count_check(port_count[1056],env.pf_vf_mux_scbd_1056.packet_count,1056);
      packet_count_check(port_count[1057],env.pf_vf_mux_scbd_1057.packet_count,1057);
      packet_count_check(port_count[1058],env.pf_vf_mux_scbd_1058.packet_count,1058);
      packet_count_check(port_count[1059],env.pf_vf_mux_scbd_1059.packet_count,1059);
      packet_count_check(port_count[1060],env.pf_vf_mux_scbd_1060.packet_count,1060);
      packet_count_check(port_count[1061],env.pf_vf_mux_scbd_1061.packet_count,1061);
      packet_count_check(port_count[1062],env.pf_vf_mux_scbd_1062.packet_count,1062);
      packet_count_check(port_count[1063],env.pf_vf_mux_scbd_1063.packet_count,1063);
      packet_count_check(port_count[1064],env.pf_vf_mux_scbd_1064.packet_count,1064);
      packet_count_check(port_count[1065],env.pf_vf_mux_scbd_1065.packet_count,1065);
      packet_count_check(port_count[1066],env.pf_vf_mux_scbd_1066.packet_count,1066);
      packet_count_check(port_count[1067],env.pf_vf_mux_scbd_1067.packet_count,1067);
      packet_count_check(port_count[1068],env.pf_vf_mux_scbd_1068.packet_count,1068);
      packet_count_check(port_count[1069],env.pf_vf_mux_scbd_1069.packet_count,1069);
      packet_count_check(port_count[1070],env.pf_vf_mux_scbd_1070.packet_count,1070);
      packet_count_check(port_count[1071],env.pf_vf_mux_scbd_1071.packet_count,1071);
      packet_count_check(port_count[1072],env.pf_vf_mux_scbd_1072.packet_count,1072);
      packet_count_check(port_count[1073],env.pf_vf_mux_scbd_1073.packet_count,1073);
      packet_count_check(port_count[1074],env.pf_vf_mux_scbd_1074.packet_count,1074);
      packet_count_check(port_count[1075],env.pf_vf_mux_scbd_1075.packet_count,1075);
      packet_count_check(port_count[1076],env.pf_vf_mux_scbd_1076.packet_count,1076);
      packet_count_check(port_count[1077],env.pf_vf_mux_scbd_1077.packet_count,1077);
      packet_count_check(port_count[1078],env.pf_vf_mux_scbd_1078.packet_count,1078);
      packet_count_check(port_count[1079],env.pf_vf_mux_scbd_1079.packet_count,1079);
      packet_count_check(port_count[1080],env.pf_vf_mux_scbd_1080.packet_count,1080);
      packet_count_check(port_count[1081],env.pf_vf_mux_scbd_1081.packet_count,1081);
      packet_count_check(port_count[1082],env.pf_vf_mux_scbd_1082.packet_count,1082);
      packet_count_check(port_count[1083],env.pf_vf_mux_scbd_1083.packet_count,1083);
      packet_count_check(port_count[1084],env.pf_vf_mux_scbd_1084.packet_count,1084);
      packet_count_check(port_count[1085],env.pf_vf_mux_scbd_1085.packet_count,1085);
      packet_count_check(port_count[1086],env.pf_vf_mux_scbd_1086.packet_count,1086);
      packet_count_check(port_count[1087],env.pf_vf_mux_scbd_1087.packet_count,1087);
      packet_count_check(port_count[1088],env.pf_vf_mux_scbd_1088.packet_count,1088);
      packet_count_check(port_count[1089],env.pf_vf_mux_scbd_1089.packet_count,1089);
      packet_count_check(port_count[1090],env.pf_vf_mux_scbd_1090.packet_count,1090);
      packet_count_check(port_count[1091],env.pf_vf_mux_scbd_1091.packet_count,1091);
      packet_count_check(port_count[1092],env.pf_vf_mux_scbd_1092.packet_count,1092);
      packet_count_check(port_count[1093],env.pf_vf_mux_scbd_1093.packet_count,1093);
      packet_count_check(port_count[1094],env.pf_vf_mux_scbd_1094.packet_count,1094);
      packet_count_check(port_count[1095],env.pf_vf_mux_scbd_1095.packet_count,1095);
      packet_count_check(port_count[1096],env.pf_vf_mux_scbd_1096.packet_count,1096);
      packet_count_check(port_count[1097],env.pf_vf_mux_scbd_1097.packet_count,1097);
      packet_count_check(port_count[1098],env.pf_vf_mux_scbd_1098.packet_count,1098);
      packet_count_check(port_count[1099],env.pf_vf_mux_scbd_1099.packet_count,1099);
      packet_count_check(port_count[1100],env.pf_vf_mux_scbd_1100.packet_count,1100);
      packet_count_check(port_count[1101],env.pf_vf_mux_scbd_1101.packet_count,1101);
      packet_count_check(port_count[1102],env.pf_vf_mux_scbd_1102.packet_count,1102);
      packet_count_check(port_count[1103],env.pf_vf_mux_scbd_1103.packet_count,1103);
      packet_count_check(port_count[1104],env.pf_vf_mux_scbd_1104.packet_count,1104);
      packet_count_check(port_count[1105],env.pf_vf_mux_scbd_1105.packet_count,1105);
      packet_count_check(port_count[1106],env.pf_vf_mux_scbd_1106.packet_count,1106);
      packet_count_check(port_count[1107],env.pf_vf_mux_scbd_1107.packet_count,1107);
      packet_count_check(port_count[1108],env.pf_vf_mux_scbd_1108.packet_count,1108);
      packet_count_check(port_count[1109],env.pf_vf_mux_scbd_1109.packet_count,1109);
      packet_count_check(port_count[1110],env.pf_vf_mux_scbd_1110.packet_count,1110);
      packet_count_check(port_count[1111],env.pf_vf_mux_scbd_1111.packet_count,1111);
      packet_count_check(port_count[1112],env.pf_vf_mux_scbd_1112.packet_count,1112);
      packet_count_check(port_count[1113],env.pf_vf_mux_scbd_1113.packet_count,1113);
      packet_count_check(port_count[1114],env.pf_vf_mux_scbd_1114.packet_count,1114);
      packet_count_check(port_count[1115],env.pf_vf_mux_scbd_1115.packet_count,1115);
      packet_count_check(port_count[1116],env.pf_vf_mux_scbd_1116.packet_count,1116);
      packet_count_check(port_count[1117],env.pf_vf_mux_scbd_1117.packet_count,1117);
      packet_count_check(port_count[1118],env.pf_vf_mux_scbd_1118.packet_count,1118);
      packet_count_check(port_count[1119],env.pf_vf_mux_scbd_1119.packet_count,1119);
      packet_count_check(port_count[1120],env.pf_vf_mux_scbd_1120.packet_count,1120);
      packet_count_check(port_count[1121],env.pf_vf_mux_scbd_1121.packet_count,1121);
      packet_count_check(port_count[1122],env.pf_vf_mux_scbd_1122.packet_count,1122);
      packet_count_check(port_count[1123],env.pf_vf_mux_scbd_1123.packet_count,1123);
      packet_count_check(port_count[1124],env.pf_vf_mux_scbd_1124.packet_count,1124);
      packet_count_check(port_count[1125],env.pf_vf_mux_scbd_1125.packet_count,1125);
      packet_count_check(port_count[1126],env.pf_vf_mux_scbd_1126.packet_count,1126);
      packet_count_check(port_count[1127],env.pf_vf_mux_scbd_1127.packet_count,1127);
      packet_count_check(port_count[1128],env.pf_vf_mux_scbd_1128.packet_count,1128);
      packet_count_check(port_count[1129],env.pf_vf_mux_scbd_1129.packet_count,1129);
      packet_count_check(port_count[1130],env.pf_vf_mux_scbd_1130.packet_count,1130);
      packet_count_check(port_count[1131],env.pf_vf_mux_scbd_1131.packet_count,1131);
      packet_count_check(port_count[1132],env.pf_vf_mux_scbd_1132.packet_count,1132);
      packet_count_check(port_count[1133],env.pf_vf_mux_scbd_1133.packet_count,1133);
      packet_count_check(port_count[1134],env.pf_vf_mux_scbd_1134.packet_count,1134);
      packet_count_check(port_count[1135],env.pf_vf_mux_scbd_1135.packet_count,1135);
      packet_count_check(port_count[1136],env.pf_vf_mux_scbd_1136.packet_count,1136);
      packet_count_check(port_count[1137],env.pf_vf_mux_scbd_1137.packet_count,1137);
      packet_count_check(port_count[1138],env.pf_vf_mux_scbd_1138.packet_count,1138);
      packet_count_check(port_count[1139],env.pf_vf_mux_scbd_1139.packet_count,1139);
      packet_count_check(port_count[1140],env.pf_vf_mux_scbd_1140.packet_count,1140);
      packet_count_check(port_count[1141],env.pf_vf_mux_scbd_1141.packet_count,1141);
      packet_count_check(port_count[1142],env.pf_vf_mux_scbd_1142.packet_count,1142);
      packet_count_check(port_count[1143],env.pf_vf_mux_scbd_1143.packet_count,1143);
      packet_count_check(port_count[1144],env.pf_vf_mux_scbd_1144.packet_count,1144);
      packet_count_check(port_count[1145],env.pf_vf_mux_scbd_1145.packet_count,1145);
      packet_count_check(port_count[1146],env.pf_vf_mux_scbd_1146.packet_count,1146);
      packet_count_check(port_count[1147],env.pf_vf_mux_scbd_1147.packet_count,1147);
      packet_count_check(port_count[1148],env.pf_vf_mux_scbd_1148.packet_count,1148);
      packet_count_check(port_count[1149],env.pf_vf_mux_scbd_1149.packet_count,1149);
      packet_count_check(port_count[1150],env.pf_vf_mux_scbd_1150.packet_count,1150);
      packet_count_check(port_count[1151],env.pf_vf_mux_scbd_1151.packet_count,1151);
      packet_count_check(port_count[1152],env.pf_vf_mux_scbd_1152.packet_count,1152);
      packet_count_check(port_count[1153],env.pf_vf_mux_scbd_1153.packet_count,1153);
      packet_count_check(port_count[1154],env.pf_vf_mux_scbd_1154.packet_count,1154);
      packet_count_check(port_count[1155],env.pf_vf_mux_scbd_1155.packet_count,1155);
      packet_count_check(port_count[1156],env.pf_vf_mux_scbd_1156.packet_count,1156);
      packet_count_check(port_count[1157],env.pf_vf_mux_scbd_1157.packet_count,1157);
      packet_count_check(port_count[1158],env.pf_vf_mux_scbd_1158.packet_count,1158);
      packet_count_check(port_count[1159],env.pf_vf_mux_scbd_1159.packet_count,1159);
      packet_count_check(port_count[1160],env.pf_vf_mux_scbd_1160.packet_count,1160);
      packet_count_check(port_count[1161],env.pf_vf_mux_scbd_1161.packet_count,1161);
      packet_count_check(port_count[1162],env.pf_vf_mux_scbd_1162.packet_count,1162);
      packet_count_check(port_count[1163],env.pf_vf_mux_scbd_1163.packet_count,1163);
      packet_count_check(port_count[1164],env.pf_vf_mux_scbd_1164.packet_count,1164);
      packet_count_check(port_count[1165],env.pf_vf_mux_scbd_1165.packet_count,1165);
      packet_count_check(port_count[1166],env.pf_vf_mux_scbd_1166.packet_count,1166);
      packet_count_check(port_count[1167],env.pf_vf_mux_scbd_1167.packet_count,1167);
      packet_count_check(port_count[1168],env.pf_vf_mux_scbd_1168.packet_count,1168);
      packet_count_check(port_count[1169],env.pf_vf_mux_scbd_1169.packet_count,1169);
      packet_count_check(port_count[1170],env.pf_vf_mux_scbd_1170.packet_count,1170);
      packet_count_check(port_count[1171],env.pf_vf_mux_scbd_1171.packet_count,1171);
      packet_count_check(port_count[1172],env.pf_vf_mux_scbd_1172.packet_count,1172);
      packet_count_check(port_count[1173],env.pf_vf_mux_scbd_1173.packet_count,1173);
      packet_count_check(port_count[1174],env.pf_vf_mux_scbd_1174.packet_count,1174);
      packet_count_check(port_count[1175],env.pf_vf_mux_scbd_1175.packet_count,1175);
      packet_count_check(port_count[1176],env.pf_vf_mux_scbd_1176.packet_count,1176);
      packet_count_check(port_count[1177],env.pf_vf_mux_scbd_1177.packet_count,1177);
      packet_count_check(port_count[1178],env.pf_vf_mux_scbd_1178.packet_count,1178);
      packet_count_check(port_count[1179],env.pf_vf_mux_scbd_1179.packet_count,1179);
      packet_count_check(port_count[1180],env.pf_vf_mux_scbd_1180.packet_count,1180);
      packet_count_check(port_count[1181],env.pf_vf_mux_scbd_1181.packet_count,1181);
      packet_count_check(port_count[1182],env.pf_vf_mux_scbd_1182.packet_count,1182);
      packet_count_check(port_count[1183],env.pf_vf_mux_scbd_1183.packet_count,1183);
      packet_count_check(port_count[1184],env.pf_vf_mux_scbd_1184.packet_count,1184);
      packet_count_check(port_count[1185],env.pf_vf_mux_scbd_1185.packet_count,1185);
      packet_count_check(port_count[1186],env.pf_vf_mux_scbd_1186.packet_count,1186);
      packet_count_check(port_count[1187],env.pf_vf_mux_scbd_1187.packet_count,1187);
      packet_count_check(port_count[1188],env.pf_vf_mux_scbd_1188.packet_count,1188);
      packet_count_check(port_count[1189],env.pf_vf_mux_scbd_1189.packet_count,1189);
      packet_count_check(port_count[1190],env.pf_vf_mux_scbd_1190.packet_count,1190);
      packet_count_check(port_count[1191],env.pf_vf_mux_scbd_1191.packet_count,1191);
      packet_count_check(port_count[1192],env.pf_vf_mux_scbd_1192.packet_count,1192);
      packet_count_check(port_count[1193],env.pf_vf_mux_scbd_1193.packet_count,1193);
      packet_count_check(port_count[1194],env.pf_vf_mux_scbd_1194.packet_count,1194);
      packet_count_check(port_count[1195],env.pf_vf_mux_scbd_1195.packet_count,1195);
      packet_count_check(port_count[1196],env.pf_vf_mux_scbd_1196.packet_count,1196);
      packet_count_check(port_count[1197],env.pf_vf_mux_scbd_1197.packet_count,1197);
      packet_count_check(port_count[1198],env.pf_vf_mux_scbd_1198.packet_count,1198);
      packet_count_check(port_count[1199],env.pf_vf_mux_scbd_1199.packet_count,1199);
      packet_count_check(port_count[1200],env.pf_vf_mux_scbd_1200.packet_count,1200);
      packet_count_check(port_count[1201],env.pf_vf_mux_scbd_1201.packet_count,1201);
      packet_count_check(port_count[1202],env.pf_vf_mux_scbd_1202.packet_count,1202);
      packet_count_check(port_count[1203],env.pf_vf_mux_scbd_1203.packet_count,1203);
      packet_count_check(port_count[1204],env.pf_vf_mux_scbd_1204.packet_count,1204);
      packet_count_check(port_count[1205],env.pf_vf_mux_scbd_1205.packet_count,1205);
      packet_count_check(port_count[1206],env.pf_vf_mux_scbd_1206.packet_count,1206);
      packet_count_check(port_count[1207],env.pf_vf_mux_scbd_1207.packet_count,1207);
      packet_count_check(port_count[1208],env.pf_vf_mux_scbd_1208.packet_count,1208);
      packet_count_check(port_count[1209],env.pf_vf_mux_scbd_1209.packet_count,1209);
      packet_count_check(port_count[1210],env.pf_vf_mux_scbd_1210.packet_count,1210);
      packet_count_check(port_count[1211],env.pf_vf_mux_scbd_1211.packet_count,1211);
      packet_count_check(port_count[1212],env.pf_vf_mux_scbd_1212.packet_count,1212);
      packet_count_check(port_count[1213],env.pf_vf_mux_scbd_1213.packet_count,1213);
      packet_count_check(port_count[1214],env.pf_vf_mux_scbd_1214.packet_count,1214);
      packet_count_check(port_count[1215],env.pf_vf_mux_scbd_1215.packet_count,1215);
      packet_count_check(port_count[1216],env.pf_vf_mux_scbd_1216.packet_count,1216);
      packet_count_check(port_count[1217],env.pf_vf_mux_scbd_1217.packet_count,1217);
      packet_count_check(port_count[1218],env.pf_vf_mux_scbd_1218.packet_count,1218);
      packet_count_check(port_count[1219],env.pf_vf_mux_scbd_1219.packet_count,1219);
      packet_count_check(port_count[1220],env.pf_vf_mux_scbd_1220.packet_count,1220);
      packet_count_check(port_count[1221],env.pf_vf_mux_scbd_1221.packet_count,1221);
      packet_count_check(port_count[1222],env.pf_vf_mux_scbd_1222.packet_count,1222);
      packet_count_check(port_count[1223],env.pf_vf_mux_scbd_1223.packet_count,1223);
      packet_count_check(port_count[1224],env.pf_vf_mux_scbd_1224.packet_count,1224);
      packet_count_check(port_count[1225],env.pf_vf_mux_scbd_1225.packet_count,1225);
      packet_count_check(port_count[1226],env.pf_vf_mux_scbd_1226.packet_count,1226);
      packet_count_check(port_count[1227],env.pf_vf_mux_scbd_1227.packet_count,1227);
      packet_count_check(port_count[1228],env.pf_vf_mux_scbd_1228.packet_count,1228);
      packet_count_check(port_count[1229],env.pf_vf_mux_scbd_1229.packet_count,1229);
      packet_count_check(port_count[1230],env.pf_vf_mux_scbd_1230.packet_count,1230);
      packet_count_check(port_count[1231],env.pf_vf_mux_scbd_1231.packet_count,1231);
      packet_count_check(port_count[1232],env.pf_vf_mux_scbd_1232.packet_count,1232);
      packet_count_check(port_count[1233],env.pf_vf_mux_scbd_1233.packet_count,1233);
      packet_count_check(port_count[1234],env.pf_vf_mux_scbd_1234.packet_count,1234);
      packet_count_check(port_count[1235],env.pf_vf_mux_scbd_1235.packet_count,1235);
      packet_count_check(port_count[1236],env.pf_vf_mux_scbd_1236.packet_count,1236);
      packet_count_check(port_count[1237],env.pf_vf_mux_scbd_1237.packet_count,1237);
      packet_count_check(port_count[1238],env.pf_vf_mux_scbd_1238.packet_count,1238);
      packet_count_check(port_count[1239],env.pf_vf_mux_scbd_1239.packet_count,1239);
      packet_count_check(port_count[1240],env.pf_vf_mux_scbd_1240.packet_count,1240);
      packet_count_check(port_count[1241],env.pf_vf_mux_scbd_1241.packet_count,1241);
      packet_count_check(port_count[1242],env.pf_vf_mux_scbd_1242.packet_count,1242);
      packet_count_check(port_count[1243],env.pf_vf_mux_scbd_1243.packet_count,1243);
      packet_count_check(port_count[1244],env.pf_vf_mux_scbd_1244.packet_count,1244);
      packet_count_check(port_count[1245],env.pf_vf_mux_scbd_1245.packet_count,1245);
      packet_count_check(port_count[1246],env.pf_vf_mux_scbd_1246.packet_count,1246);
      packet_count_check(port_count[1247],env.pf_vf_mux_scbd_1247.packet_count,1247);
      packet_count_check(port_count[1248],env.pf_vf_mux_scbd_1248.packet_count,1248);
      packet_count_check(port_count[1249],env.pf_vf_mux_scbd_1249.packet_count,1249);
      packet_count_check(port_count[1250],env.pf_vf_mux_scbd_1250.packet_count,1250);
      packet_count_check(port_count[1251],env.pf_vf_mux_scbd_1251.packet_count,1251);
      packet_count_check(port_count[1252],env.pf_vf_mux_scbd_1252.packet_count,1252);
      packet_count_check(port_count[1253],env.pf_vf_mux_scbd_1253.packet_count,1253);
      packet_count_check(port_count[1254],env.pf_vf_mux_scbd_1254.packet_count,1254);
      packet_count_check(port_count[1255],env.pf_vf_mux_scbd_1255.packet_count,1255);
      packet_count_check(port_count[1256],env.pf_vf_mux_scbd_1256.packet_count,1256);
      packet_count_check(port_count[1257],env.pf_vf_mux_scbd_1257.packet_count,1257);
      packet_count_check(port_count[1258],env.pf_vf_mux_scbd_1258.packet_count,1258);
      packet_count_check(port_count[1259],env.pf_vf_mux_scbd_1259.packet_count,1259);
      packet_count_check(port_count[1260],env.pf_vf_mux_scbd_1260.packet_count,1260);
      packet_count_check(port_count[1261],env.pf_vf_mux_scbd_1261.packet_count,1261);
      packet_count_check(port_count[1262],env.pf_vf_mux_scbd_1262.packet_count,1262);
      packet_count_check(port_count[1263],env.pf_vf_mux_scbd_1263.packet_count,1263);
      packet_count_check(port_count[1264],env.pf_vf_mux_scbd_1264.packet_count,1264);
      packet_count_check(port_count[1265],env.pf_vf_mux_scbd_1265.packet_count,1265);
      packet_count_check(port_count[1266],env.pf_vf_mux_scbd_1266.packet_count,1266);
      packet_count_check(port_count[1267],env.pf_vf_mux_scbd_1267.packet_count,1267);
      packet_count_check(port_count[1268],env.pf_vf_mux_scbd_1268.packet_count,1268);
      packet_count_check(port_count[1269],env.pf_vf_mux_scbd_1269.packet_count,1269);
      packet_count_check(port_count[1270],env.pf_vf_mux_scbd_1270.packet_count,1270);
      packet_count_check(port_count[1271],env.pf_vf_mux_scbd_1271.packet_count,1271);
      packet_count_check(port_count[1272],env.pf_vf_mux_scbd_1272.packet_count,1272);
      packet_count_check(port_count[1273],env.pf_vf_mux_scbd_1273.packet_count,1273);
      packet_count_check(port_count[1274],env.pf_vf_mux_scbd_1274.packet_count,1274);
      packet_count_check(port_count[1275],env.pf_vf_mux_scbd_1275.packet_count,1275);
      packet_count_check(port_count[1276],env.pf_vf_mux_scbd_1276.packet_count,1276);
      packet_count_check(port_count[1277],env.pf_vf_mux_scbd_1277.packet_count,1277);
      packet_count_check(port_count[1278],env.pf_vf_mux_scbd_1278.packet_count,1278);
      packet_count_check(port_count[1279],env.pf_vf_mux_scbd_1279.packet_count,1279);
      packet_count_check(port_count[1280],env.pf_vf_mux_scbd_1280.packet_count,1280);
      packet_count_check(port_count[1281],env.pf_vf_mux_scbd_1281.packet_count,1281);
      packet_count_check(port_count[1282],env.pf_vf_mux_scbd_1282.packet_count,1282);
      packet_count_check(port_count[1283],env.pf_vf_mux_scbd_1283.packet_count,1283);
      packet_count_check(port_count[1284],env.pf_vf_mux_scbd_1284.packet_count,1284);
      packet_count_check(port_count[1285],env.pf_vf_mux_scbd_1285.packet_count,1285);
      packet_count_check(port_count[1286],env.pf_vf_mux_scbd_1286.packet_count,1286);
      packet_count_check(port_count[1287],env.pf_vf_mux_scbd_1287.packet_count,1287);
      packet_count_check(port_count[1288],env.pf_vf_mux_scbd_1288.packet_count,1288);
      packet_count_check(port_count[1289],env.pf_vf_mux_scbd_1289.packet_count,1289);
      packet_count_check(port_count[1290],env.pf_vf_mux_scbd_1290.packet_count,1290);
      packet_count_check(port_count[1291],env.pf_vf_mux_scbd_1291.packet_count,1291);
      packet_count_check(port_count[1292],env.pf_vf_mux_scbd_1292.packet_count,1292);
      packet_count_check(port_count[1293],env.pf_vf_mux_scbd_1293.packet_count,1293);
      packet_count_check(port_count[1294],env.pf_vf_mux_scbd_1294.packet_count,1294);
      packet_count_check(port_count[1295],env.pf_vf_mux_scbd_1295.packet_count,1295);
      packet_count_check(port_count[1296],env.pf_vf_mux_scbd_1296.packet_count,1296);
      packet_count_check(port_count[1297],env.pf_vf_mux_scbd_1297.packet_count,1297);
      packet_count_check(port_count[1298],env.pf_vf_mux_scbd_1298.packet_count,1298);
      packet_count_check(port_count[1299],env.pf_vf_mux_scbd_1299.packet_count,1299);
      packet_count_check(port_count[1300],env.pf_vf_mux_scbd_1300.packet_count,1300);
      packet_count_check(port_count[1301],env.pf_vf_mux_scbd_1301.packet_count,1301);
      packet_count_check(port_count[1302],env.pf_vf_mux_scbd_1302.packet_count,1302);
      packet_count_check(port_count[1303],env.pf_vf_mux_scbd_1303.packet_count,1303);
      packet_count_check(port_count[1304],env.pf_vf_mux_scbd_1304.packet_count,1304);
      packet_count_check(port_count[1305],env.pf_vf_mux_scbd_1305.packet_count,1305);
      packet_count_check(port_count[1306],env.pf_vf_mux_scbd_1306.packet_count,1306);
      packet_count_check(port_count[1307],env.pf_vf_mux_scbd_1307.packet_count,1307);
      packet_count_check(port_count[1308],env.pf_vf_mux_scbd_1308.packet_count,1308);
      packet_count_check(port_count[1309],env.pf_vf_mux_scbd_1309.packet_count,1309);
      packet_count_check(port_count[1310],env.pf_vf_mux_scbd_1310.packet_count,1310);
      packet_count_check(port_count[1311],env.pf_vf_mux_scbd_1311.packet_count,1311);
      packet_count_check(port_count[1312],env.pf_vf_mux_scbd_1312.packet_count,1312);
      packet_count_check(port_count[1313],env.pf_vf_mux_scbd_1313.packet_count,1313);
      packet_count_check(port_count[1314],env.pf_vf_mux_scbd_1314.packet_count,1314);
      packet_count_check(port_count[1315],env.pf_vf_mux_scbd_1315.packet_count,1315);
      packet_count_check(port_count[1316],env.pf_vf_mux_scbd_1316.packet_count,1316);
      packet_count_check(port_count[1317],env.pf_vf_mux_scbd_1317.packet_count,1317);
      packet_count_check(port_count[1318],env.pf_vf_mux_scbd_1318.packet_count,1318);
      packet_count_check(port_count[1319],env.pf_vf_mux_scbd_1319.packet_count,1319);
      packet_count_check(port_count[1320],env.pf_vf_mux_scbd_1320.packet_count,1320);
      packet_count_check(port_count[1321],env.pf_vf_mux_scbd_1321.packet_count,1321);
      packet_count_check(port_count[1322],env.pf_vf_mux_scbd_1322.packet_count,1322);
      packet_count_check(port_count[1323],env.pf_vf_mux_scbd_1323.packet_count,1323);
      packet_count_check(port_count[1324],env.pf_vf_mux_scbd_1324.packet_count,1324);
      packet_count_check(port_count[1325],env.pf_vf_mux_scbd_1325.packet_count,1325);
      packet_count_check(port_count[1326],env.pf_vf_mux_scbd_1326.packet_count,1326);
      packet_count_check(port_count[1327],env.pf_vf_mux_scbd_1327.packet_count,1327);
      packet_count_check(port_count[1328],env.pf_vf_mux_scbd_1328.packet_count,1328);
      packet_count_check(port_count[1329],env.pf_vf_mux_scbd_1329.packet_count,1329);
      packet_count_check(port_count[1330],env.pf_vf_mux_scbd_1330.packet_count,1330);
      packet_count_check(port_count[1331],env.pf_vf_mux_scbd_1331.packet_count,1331);
      packet_count_check(port_count[1332],env.pf_vf_mux_scbd_1332.packet_count,1332);
      packet_count_check(port_count[1333],env.pf_vf_mux_scbd_1333.packet_count,1333);
      packet_count_check(port_count[1334],env.pf_vf_mux_scbd_1334.packet_count,1334);
      packet_count_check(port_count[1335],env.pf_vf_mux_scbd_1335.packet_count,1335);
      packet_count_check(port_count[1336],env.pf_vf_mux_scbd_1336.packet_count,1336);
      packet_count_check(port_count[1337],env.pf_vf_mux_scbd_1337.packet_count,1337);
      packet_count_check(port_count[1338],env.pf_vf_mux_scbd_1338.packet_count,1338);
      packet_count_check(port_count[1339],env.pf_vf_mux_scbd_1339.packet_count,1339);
      packet_count_check(port_count[1340],env.pf_vf_mux_scbd_1340.packet_count,1340);
      packet_count_check(port_count[1341],env.pf_vf_mux_scbd_1341.packet_count,1341);
      packet_count_check(port_count[1342],env.pf_vf_mux_scbd_1342.packet_count,1342);
      packet_count_check(port_count[1343],env.pf_vf_mux_scbd_1343.packet_count,1343);
      packet_count_check(port_count[1344],env.pf_vf_mux_scbd_1344.packet_count,1344);
      packet_count_check(port_count[1345],env.pf_vf_mux_scbd_1345.packet_count,1345);
      packet_count_check(port_count[1346],env.pf_vf_mux_scbd_1346.packet_count,1346);
      packet_count_check(port_count[1347],env.pf_vf_mux_scbd_1347.packet_count,1347);
      packet_count_check(port_count[1348],env.pf_vf_mux_scbd_1348.packet_count,1348);
      packet_count_check(port_count[1349],env.pf_vf_mux_scbd_1349.packet_count,1349);
      packet_count_check(port_count[1350],env.pf_vf_mux_scbd_1350.packet_count,1350);
      packet_count_check(port_count[1351],env.pf_vf_mux_scbd_1351.packet_count,1351);
      packet_count_check(port_count[1352],env.pf_vf_mux_scbd_1352.packet_count,1352);
      packet_count_check(port_count[1353],env.pf_vf_mux_scbd_1353.packet_count,1353);
      packet_count_check(port_count[1354],env.pf_vf_mux_scbd_1354.packet_count,1354);
      packet_count_check(port_count[1355],env.pf_vf_mux_scbd_1355.packet_count,1355);
      packet_count_check(port_count[1356],env.pf_vf_mux_scbd_1356.packet_count,1356);
      packet_count_check(port_count[1357],env.pf_vf_mux_scbd_1357.packet_count,1357);
      packet_count_check(port_count[1358],env.pf_vf_mux_scbd_1358.packet_count,1358);
      packet_count_check(port_count[1359],env.pf_vf_mux_scbd_1359.packet_count,1359);
      packet_count_check(port_count[1360],env.pf_vf_mux_scbd_1360.packet_count,1360);
      packet_count_check(port_count[1361],env.pf_vf_mux_scbd_1361.packet_count,1361);
      packet_count_check(port_count[1362],env.pf_vf_mux_scbd_1362.packet_count,1362);
      packet_count_check(port_count[1363],env.pf_vf_mux_scbd_1363.packet_count,1363);
      packet_count_check(port_count[1364],env.pf_vf_mux_scbd_1364.packet_count,1364);
      packet_count_check(port_count[1365],env.pf_vf_mux_scbd_1365.packet_count,1365);
      packet_count_check(port_count[1366],env.pf_vf_mux_scbd_1366.packet_count,1366);
      packet_count_check(port_count[1367],env.pf_vf_mux_scbd_1367.packet_count,1367);
      packet_count_check(port_count[1368],env.pf_vf_mux_scbd_1368.packet_count,1368);
      packet_count_check(port_count[1369],env.pf_vf_mux_scbd_1369.packet_count,1369);
      packet_count_check(port_count[1370],env.pf_vf_mux_scbd_1370.packet_count,1370);
      packet_count_check(port_count[1371],env.pf_vf_mux_scbd_1371.packet_count,1371);
      packet_count_check(port_count[1372],env.pf_vf_mux_scbd_1372.packet_count,1372);
      packet_count_check(port_count[1373],env.pf_vf_mux_scbd_1373.packet_count,1373);
      packet_count_check(port_count[1374],env.pf_vf_mux_scbd_1374.packet_count,1374);
      packet_count_check(port_count[1375],env.pf_vf_mux_scbd_1375.packet_count,1375);
      packet_count_check(port_count[1376],env.pf_vf_mux_scbd_1376.packet_count,1376);
      packet_count_check(port_count[1377],env.pf_vf_mux_scbd_1377.packet_count,1377);
      packet_count_check(port_count[1378],env.pf_vf_mux_scbd_1378.packet_count,1378);
      packet_count_check(port_count[1379],env.pf_vf_mux_scbd_1379.packet_count,1379);
      packet_count_check(port_count[1380],env.pf_vf_mux_scbd_1380.packet_count,1380);
      packet_count_check(port_count[1381],env.pf_vf_mux_scbd_1381.packet_count,1381);
      packet_count_check(port_count[1382],env.pf_vf_mux_scbd_1382.packet_count,1382);
      packet_count_check(port_count[1383],env.pf_vf_mux_scbd_1383.packet_count,1383);
      packet_count_check(port_count[1384],env.pf_vf_mux_scbd_1384.packet_count,1384);
      packet_count_check(port_count[1385],env.pf_vf_mux_scbd_1385.packet_count,1385);
      packet_count_check(port_count[1386],env.pf_vf_mux_scbd_1386.packet_count,1386);
      packet_count_check(port_count[1387],env.pf_vf_mux_scbd_1387.packet_count,1387);
      packet_count_check(port_count[1388],env.pf_vf_mux_scbd_1388.packet_count,1388);
      packet_count_check(port_count[1389],env.pf_vf_mux_scbd_1389.packet_count,1389);
      packet_count_check(port_count[1390],env.pf_vf_mux_scbd_1390.packet_count,1390);
      packet_count_check(port_count[1391],env.pf_vf_mux_scbd_1391.packet_count,1391);
      packet_count_check(port_count[1392],env.pf_vf_mux_scbd_1392.packet_count,1392);
      packet_count_check(port_count[1393],env.pf_vf_mux_scbd_1393.packet_count,1393);
      packet_count_check(port_count[1394],env.pf_vf_mux_scbd_1394.packet_count,1394);
      packet_count_check(port_count[1395],env.pf_vf_mux_scbd_1395.packet_count,1395);
      packet_count_check(port_count[1396],env.pf_vf_mux_scbd_1396.packet_count,1396);
      packet_count_check(port_count[1397],env.pf_vf_mux_scbd_1397.packet_count,1397);
      packet_count_check(port_count[1398],env.pf_vf_mux_scbd_1398.packet_count,1398);
      packet_count_check(port_count[1399],env.pf_vf_mux_scbd_1399.packet_count,1399);
      packet_count_check(port_count[1400],env.pf_vf_mux_scbd_1400.packet_count,1400);
      packet_count_check(port_count[1401],env.pf_vf_mux_scbd_1401.packet_count,1401);
      packet_count_check(port_count[1402],env.pf_vf_mux_scbd_1402.packet_count,1402);
      packet_count_check(port_count[1403],env.pf_vf_mux_scbd_1403.packet_count,1403);
      packet_count_check(port_count[1404],env.pf_vf_mux_scbd_1404.packet_count,1404);
      packet_count_check(port_count[1405],env.pf_vf_mux_scbd_1405.packet_count,1405);
      packet_count_check(port_count[1406],env.pf_vf_mux_scbd_1406.packet_count,1406);
      packet_count_check(port_count[1407],env.pf_vf_mux_scbd_1407.packet_count,1407);
      packet_count_check(port_count[1408],env.pf_vf_mux_scbd_1408.packet_count,1408);
      packet_count_check(port_count[1409],env.pf_vf_mux_scbd_1409.packet_count,1409);
      packet_count_check(port_count[1410],env.pf_vf_mux_scbd_1410.packet_count,1410);
      packet_count_check(port_count[1411],env.pf_vf_mux_scbd_1411.packet_count,1411);
      packet_count_check(port_count[1412],env.pf_vf_mux_scbd_1412.packet_count,1412);
      packet_count_check(port_count[1413],env.pf_vf_mux_scbd_1413.packet_count,1413);
      packet_count_check(port_count[1414],env.pf_vf_mux_scbd_1414.packet_count,1414);
      packet_count_check(port_count[1415],env.pf_vf_mux_scbd_1415.packet_count,1415);
      packet_count_check(port_count[1416],env.pf_vf_mux_scbd_1416.packet_count,1416);
      packet_count_check(port_count[1417],env.pf_vf_mux_scbd_1417.packet_count,1417);
      packet_count_check(port_count[1418],env.pf_vf_mux_scbd_1418.packet_count,1418);
      packet_count_check(port_count[1419],env.pf_vf_mux_scbd_1419.packet_count,1419);
      packet_count_check(port_count[1420],env.pf_vf_mux_scbd_1420.packet_count,1420);
      packet_count_check(port_count[1421],env.pf_vf_mux_scbd_1421.packet_count,1421);
      packet_count_check(port_count[1422],env.pf_vf_mux_scbd_1422.packet_count,1422);
      packet_count_check(port_count[1423],env.pf_vf_mux_scbd_1423.packet_count,1423);
      packet_count_check(port_count[1424],env.pf_vf_mux_scbd_1424.packet_count,1424);
      packet_count_check(port_count[1425],env.pf_vf_mux_scbd_1425.packet_count,1425);
      packet_count_check(port_count[1426],env.pf_vf_mux_scbd_1426.packet_count,1426);
      packet_count_check(port_count[1427],env.pf_vf_mux_scbd_1427.packet_count,1427);
      packet_count_check(port_count[1428],env.pf_vf_mux_scbd_1428.packet_count,1428);
      packet_count_check(port_count[1429],env.pf_vf_mux_scbd_1429.packet_count,1429);
      packet_count_check(port_count[1430],env.pf_vf_mux_scbd_1430.packet_count,1430);
      packet_count_check(port_count[1431],env.pf_vf_mux_scbd_1431.packet_count,1431);
      packet_count_check(port_count[1432],env.pf_vf_mux_scbd_1432.packet_count,1432);
      packet_count_check(port_count[1433],env.pf_vf_mux_scbd_1433.packet_count,1433);
      packet_count_check(port_count[1434],env.pf_vf_mux_scbd_1434.packet_count,1434);
      packet_count_check(port_count[1435],env.pf_vf_mux_scbd_1435.packet_count,1435);
      packet_count_check(port_count[1436],env.pf_vf_mux_scbd_1436.packet_count,1436);
      packet_count_check(port_count[1437],env.pf_vf_mux_scbd_1437.packet_count,1437);
      packet_count_check(port_count[1438],env.pf_vf_mux_scbd_1438.packet_count,1438);
      packet_count_check(port_count[1439],env.pf_vf_mux_scbd_1439.packet_count,1439);
      packet_count_check(port_count[1440],env.pf_vf_mux_scbd_1440.packet_count,1440);
      packet_count_check(port_count[1441],env.pf_vf_mux_scbd_1441.packet_count,1441);
      packet_count_check(port_count[1442],env.pf_vf_mux_scbd_1442.packet_count,1442);
      packet_count_check(port_count[1443],env.pf_vf_mux_scbd_1443.packet_count,1443);
      packet_count_check(port_count[1444],env.pf_vf_mux_scbd_1444.packet_count,1444);
      packet_count_check(port_count[1445],env.pf_vf_mux_scbd_1445.packet_count,1445);
      packet_count_check(port_count[1446],env.pf_vf_mux_scbd_1446.packet_count,1446);
      packet_count_check(port_count[1447],env.pf_vf_mux_scbd_1447.packet_count,1447);
      packet_count_check(port_count[1448],env.pf_vf_mux_scbd_1448.packet_count,1448);
      packet_count_check(port_count[1449],env.pf_vf_mux_scbd_1449.packet_count,1449);
      packet_count_check(port_count[1450],env.pf_vf_mux_scbd_1450.packet_count,1450);
      packet_count_check(port_count[1451],env.pf_vf_mux_scbd_1451.packet_count,1451);
      packet_count_check(port_count[1452],env.pf_vf_mux_scbd_1452.packet_count,1452);
      packet_count_check(port_count[1453],env.pf_vf_mux_scbd_1453.packet_count,1453);
      packet_count_check(port_count[1454],env.pf_vf_mux_scbd_1454.packet_count,1454);
      packet_count_check(port_count[1455],env.pf_vf_mux_scbd_1455.packet_count,1455);
      packet_count_check(port_count[1456],env.pf_vf_mux_scbd_1456.packet_count,1456);
      packet_count_check(port_count[1457],env.pf_vf_mux_scbd_1457.packet_count,1457);
      packet_count_check(port_count[1458],env.pf_vf_mux_scbd_1458.packet_count,1458);
      packet_count_check(port_count[1459],env.pf_vf_mux_scbd_1459.packet_count,1459);
      packet_count_check(port_count[1460],env.pf_vf_mux_scbd_1460.packet_count,1460);
      packet_count_check(port_count[1461],env.pf_vf_mux_scbd_1461.packet_count,1461);
      packet_count_check(port_count[1462],env.pf_vf_mux_scbd_1462.packet_count,1462);
      packet_count_check(port_count[1463],env.pf_vf_mux_scbd_1463.packet_count,1463);
      packet_count_check(port_count[1464],env.pf_vf_mux_scbd_1464.packet_count,1464);
      packet_count_check(port_count[1465],env.pf_vf_mux_scbd_1465.packet_count,1465);
      packet_count_check(port_count[1466],env.pf_vf_mux_scbd_1466.packet_count,1466);
      packet_count_check(port_count[1467],env.pf_vf_mux_scbd_1467.packet_count,1467);
      packet_count_check(port_count[1468],env.pf_vf_mux_scbd_1468.packet_count,1468);
      packet_count_check(port_count[1469],env.pf_vf_mux_scbd_1469.packet_count,1469);
      packet_count_check(port_count[1470],env.pf_vf_mux_scbd_1470.packet_count,1470);
      packet_count_check(port_count[1471],env.pf_vf_mux_scbd_1471.packet_count,1471);
      packet_count_check(port_count[1472],env.pf_vf_mux_scbd_1472.packet_count,1472);
      packet_count_check(port_count[1473],env.pf_vf_mux_scbd_1473.packet_count,1473);
      packet_count_check(port_count[1474],env.pf_vf_mux_scbd_1474.packet_count,1474);
      packet_count_check(port_count[1475],env.pf_vf_mux_scbd_1475.packet_count,1475);
      packet_count_check(port_count[1476],env.pf_vf_mux_scbd_1476.packet_count,1476);
      packet_count_check(port_count[1477],env.pf_vf_mux_scbd_1477.packet_count,1477);
      packet_count_check(port_count[1478],env.pf_vf_mux_scbd_1478.packet_count,1478);
      packet_count_check(port_count[1479],env.pf_vf_mux_scbd_1479.packet_count,1479);
      packet_count_check(port_count[1480],env.pf_vf_mux_scbd_1480.packet_count,1480);
      packet_count_check(port_count[1481],env.pf_vf_mux_scbd_1481.packet_count,1481);
      packet_count_check(port_count[1482],env.pf_vf_mux_scbd_1482.packet_count,1482);
      packet_count_check(port_count[1483],env.pf_vf_mux_scbd_1483.packet_count,1483);
      packet_count_check(port_count[1484],env.pf_vf_mux_scbd_1484.packet_count,1484);
      packet_count_check(port_count[1485],env.pf_vf_mux_scbd_1485.packet_count,1485);
      packet_count_check(port_count[1486],env.pf_vf_mux_scbd_1486.packet_count,1486);
      packet_count_check(port_count[1487],env.pf_vf_mux_scbd_1487.packet_count,1487);
      packet_count_check(port_count[1488],env.pf_vf_mux_scbd_1488.packet_count,1488);
      packet_count_check(port_count[1489],env.pf_vf_mux_scbd_1489.packet_count,1489);
      packet_count_check(port_count[1490],env.pf_vf_mux_scbd_1490.packet_count,1490);
      packet_count_check(port_count[1491],env.pf_vf_mux_scbd_1491.packet_count,1491);
      packet_count_check(port_count[1492],env.pf_vf_mux_scbd_1492.packet_count,1492);
      packet_count_check(port_count[1493],env.pf_vf_mux_scbd_1493.packet_count,1493);
      packet_count_check(port_count[1494],env.pf_vf_mux_scbd_1494.packet_count,1494);
      packet_count_check(port_count[1495],env.pf_vf_mux_scbd_1495.packet_count,1495);
      packet_count_check(port_count[1496],env.pf_vf_mux_scbd_1496.packet_count,1496);
      packet_count_check(port_count[1497],env.pf_vf_mux_scbd_1497.packet_count,1497);
      packet_count_check(port_count[1498],env.pf_vf_mux_scbd_1498.packet_count,1498);
      packet_count_check(port_count[1499],env.pf_vf_mux_scbd_1499.packet_count,1499);
      packet_count_check(port_count[1500],env.pf_vf_mux_scbd_1500.packet_count,1500);
      packet_count_check(port_count[1501],env.pf_vf_mux_scbd_1501.packet_count,1501);
      packet_count_check(port_count[1502],env.pf_vf_mux_scbd_1502.packet_count,1502);
      packet_count_check(port_count[1503],env.pf_vf_mux_scbd_1503.packet_count,1503);
      packet_count_check(port_count[1504],env.pf_vf_mux_scbd_1504.packet_count,1504);
      packet_count_check(port_count[1505],env.pf_vf_mux_scbd_1505.packet_count,1505);
      packet_count_check(port_count[1506],env.pf_vf_mux_scbd_1506.packet_count,1506);
      packet_count_check(port_count[1507],env.pf_vf_mux_scbd_1507.packet_count,1507);
      packet_count_check(port_count[1508],env.pf_vf_mux_scbd_1508.packet_count,1508);
      packet_count_check(port_count[1509],env.pf_vf_mux_scbd_1509.packet_count,1509);
      packet_count_check(port_count[1510],env.pf_vf_mux_scbd_1510.packet_count,1510);
      packet_count_check(port_count[1511],env.pf_vf_mux_scbd_1511.packet_count,1511);
      packet_count_check(port_count[1512],env.pf_vf_mux_scbd_1512.packet_count,1512);
      packet_count_check(port_count[1513],env.pf_vf_mux_scbd_1513.packet_count,1513);
      packet_count_check(port_count[1514],env.pf_vf_mux_scbd_1514.packet_count,1514);
      packet_count_check(port_count[1515],env.pf_vf_mux_scbd_1515.packet_count,1515);
      packet_count_check(port_count[1516],env.pf_vf_mux_scbd_1516.packet_count,1516);
      packet_count_check(port_count[1517],env.pf_vf_mux_scbd_1517.packet_count,1517);
      packet_count_check(port_count[1518],env.pf_vf_mux_scbd_1518.packet_count,1518);
      packet_count_check(port_count[1519],env.pf_vf_mux_scbd_1519.packet_count,1519);
      packet_count_check(port_count[1520],env.pf_vf_mux_scbd_1520.packet_count,1520);
      packet_count_check(port_count[1521],env.pf_vf_mux_scbd_1521.packet_count,1521);
      packet_count_check(port_count[1522],env.pf_vf_mux_scbd_1522.packet_count,1522);
      packet_count_check(port_count[1523],env.pf_vf_mux_scbd_1523.packet_count,1523);
      packet_count_check(port_count[1524],env.pf_vf_mux_scbd_1524.packet_count,1524);
      packet_count_check(port_count[1525],env.pf_vf_mux_scbd_1525.packet_count,1525);
      packet_count_check(port_count[1526],env.pf_vf_mux_scbd_1526.packet_count,1526);
      packet_count_check(port_count[1527],env.pf_vf_mux_scbd_1527.packet_count,1527);
      packet_count_check(port_count[1528],env.pf_vf_mux_scbd_1528.packet_count,1528);
      packet_count_check(port_count[1529],env.pf_vf_mux_scbd_1529.packet_count,1529);
      packet_count_check(port_count[1530],env.pf_vf_mux_scbd_1530.packet_count,1530);
      packet_count_check(port_count[1531],env.pf_vf_mux_scbd_1531.packet_count,1531);
      packet_count_check(port_count[1532],env.pf_vf_mux_scbd_1532.packet_count,1532);
      packet_count_check(port_count[1533],env.pf_vf_mux_scbd_1533.packet_count,1533);
      packet_count_check(port_count[1534],env.pf_vf_mux_scbd_1534.packet_count,1534);
      packet_count_check(port_count[1535],env.pf_vf_mux_scbd_1535.packet_count,1535);
      packet_count_check(port_count[1536],env.pf_vf_mux_scbd_1536.packet_count,1536);
      packet_count_check(port_count[1537],env.pf_vf_mux_scbd_1537.packet_count,1537);
      packet_count_check(port_count[1538],env.pf_vf_mux_scbd_1538.packet_count,1538);
      packet_count_check(port_count[1539],env.pf_vf_mux_scbd_1539.packet_count,1539);
      packet_count_check(port_count[1540],env.pf_vf_mux_scbd_1540.packet_count,1540);
      packet_count_check(port_count[1541],env.pf_vf_mux_scbd_1541.packet_count,1541);
      packet_count_check(port_count[1542],env.pf_vf_mux_scbd_1542.packet_count,1542);
      packet_count_check(port_count[1543],env.pf_vf_mux_scbd_1543.packet_count,1543);
      packet_count_check(port_count[1544],env.pf_vf_mux_scbd_1544.packet_count,1544);
      packet_count_check(port_count[1545],env.pf_vf_mux_scbd_1545.packet_count,1545);
      packet_count_check(port_count[1546],env.pf_vf_mux_scbd_1546.packet_count,1546);
      packet_count_check(port_count[1547],env.pf_vf_mux_scbd_1547.packet_count,1547);
      packet_count_check(port_count[1548],env.pf_vf_mux_scbd_1548.packet_count,1548);
      packet_count_check(port_count[1549],env.pf_vf_mux_scbd_1549.packet_count,1549);
      packet_count_check(port_count[1550],env.pf_vf_mux_scbd_1550.packet_count,1550);
      packet_count_check(port_count[1551],env.pf_vf_mux_scbd_1551.packet_count,1551);
      packet_count_check(port_count[1552],env.pf_vf_mux_scbd_1552.packet_count,1552);
      packet_count_check(port_count[1553],env.pf_vf_mux_scbd_1553.packet_count,1553);
      packet_count_check(port_count[1554],env.pf_vf_mux_scbd_1554.packet_count,1554);
      packet_count_check(port_count[1555],env.pf_vf_mux_scbd_1555.packet_count,1555);
      packet_count_check(port_count[1556],env.pf_vf_mux_scbd_1556.packet_count,1556);
      packet_count_check(port_count[1557],env.pf_vf_mux_scbd_1557.packet_count,1557);
      packet_count_check(port_count[1558],env.pf_vf_mux_scbd_1558.packet_count,1558);
      packet_count_check(port_count[1559],env.pf_vf_mux_scbd_1559.packet_count,1559);
      packet_count_check(port_count[1560],env.pf_vf_mux_scbd_1560.packet_count,1560);
      packet_count_check(port_count[1561],env.pf_vf_mux_scbd_1561.packet_count,1561);
      packet_count_check(port_count[1562],env.pf_vf_mux_scbd_1562.packet_count,1562);
      packet_count_check(port_count[1563],env.pf_vf_mux_scbd_1563.packet_count,1563);
      packet_count_check(port_count[1564],env.pf_vf_mux_scbd_1564.packet_count,1564);
      packet_count_check(port_count[1565],env.pf_vf_mux_scbd_1565.packet_count,1565);
      packet_count_check(port_count[1566],env.pf_vf_mux_scbd_1566.packet_count,1566);
      packet_count_check(port_count[1567],env.pf_vf_mux_scbd_1567.packet_count,1567);
      packet_count_check(port_count[1568],env.pf_vf_mux_scbd_1568.packet_count,1568);
      packet_count_check(port_count[1569],env.pf_vf_mux_scbd_1569.packet_count,1569);
      packet_count_check(port_count[1570],env.pf_vf_mux_scbd_1570.packet_count,1570);
      packet_count_check(port_count[1571],env.pf_vf_mux_scbd_1571.packet_count,1571);
      packet_count_check(port_count[1572],env.pf_vf_mux_scbd_1572.packet_count,1572);
      packet_count_check(port_count[1573],env.pf_vf_mux_scbd_1573.packet_count,1573);
      packet_count_check(port_count[1574],env.pf_vf_mux_scbd_1574.packet_count,1574);
      packet_count_check(port_count[1575],env.pf_vf_mux_scbd_1575.packet_count,1575);
      packet_count_check(port_count[1576],env.pf_vf_mux_scbd_1576.packet_count,1576);
      packet_count_check(port_count[1577],env.pf_vf_mux_scbd_1577.packet_count,1577);
      packet_count_check(port_count[1578],env.pf_vf_mux_scbd_1578.packet_count,1578);
      packet_count_check(port_count[1579],env.pf_vf_mux_scbd_1579.packet_count,1579);
      packet_count_check(port_count[1580],env.pf_vf_mux_scbd_1580.packet_count,1580);
      packet_count_check(port_count[1581],env.pf_vf_mux_scbd_1581.packet_count,1581);
      packet_count_check(port_count[1582],env.pf_vf_mux_scbd_1582.packet_count,1582);
      packet_count_check(port_count[1583],env.pf_vf_mux_scbd_1583.packet_count,1583);
      packet_count_check(port_count[1584],env.pf_vf_mux_scbd_1584.packet_count,1584);
      packet_count_check(port_count[1585],env.pf_vf_mux_scbd_1585.packet_count,1585);
      packet_count_check(port_count[1586],env.pf_vf_mux_scbd_1586.packet_count,1586);
      packet_count_check(port_count[1587],env.pf_vf_mux_scbd_1587.packet_count,1587);
      packet_count_check(port_count[1588],env.pf_vf_mux_scbd_1588.packet_count,1588);
      packet_count_check(port_count[1589],env.pf_vf_mux_scbd_1589.packet_count,1589);
      packet_count_check(port_count[1590],env.pf_vf_mux_scbd_1590.packet_count,1590);
      packet_count_check(port_count[1591],env.pf_vf_mux_scbd_1591.packet_count,1591);
      packet_count_check(port_count[1592],env.pf_vf_mux_scbd_1592.packet_count,1592);
      packet_count_check(port_count[1593],env.pf_vf_mux_scbd_1593.packet_count,1593);
      packet_count_check(port_count[1594],env.pf_vf_mux_scbd_1594.packet_count,1594);
      packet_count_check(port_count[1595],env.pf_vf_mux_scbd_1595.packet_count,1595);
      packet_count_check(port_count[1596],env.pf_vf_mux_scbd_1596.packet_count,1596);
      packet_count_check(port_count[1597],env.pf_vf_mux_scbd_1597.packet_count,1597);
      packet_count_check(port_count[1598],env.pf_vf_mux_scbd_1598.packet_count,1598);
      packet_count_check(port_count[1599],env.pf_vf_mux_scbd_1599.packet_count,1599);
      packet_count_check(port_count[1600],env.pf_vf_mux_scbd_1600.packet_count,1600);
      packet_count_check(port_count[1601],env.pf_vf_mux_scbd_1601.packet_count,1601);
      packet_count_check(port_count[1602],env.pf_vf_mux_scbd_1602.packet_count,1602);
      packet_count_check(port_count[1603],env.pf_vf_mux_scbd_1603.packet_count,1603);
      packet_count_check(port_count[1604],env.pf_vf_mux_scbd_1604.packet_count,1604);
      packet_count_check(port_count[1605],env.pf_vf_mux_scbd_1605.packet_count,1605);
      packet_count_check(port_count[1606],env.pf_vf_mux_scbd_1606.packet_count,1606);
      packet_count_check(port_count[1607],env.pf_vf_mux_scbd_1607.packet_count,1607);
      packet_count_check(port_count[1608],env.pf_vf_mux_scbd_1608.packet_count,1608);
      packet_count_check(port_count[1609],env.pf_vf_mux_scbd_1609.packet_count,1609);
      packet_count_check(port_count[1610],env.pf_vf_mux_scbd_1610.packet_count,1610);
      packet_count_check(port_count[1611],env.pf_vf_mux_scbd_1611.packet_count,1611);
      packet_count_check(port_count[1612],env.pf_vf_mux_scbd_1612.packet_count,1612);
      packet_count_check(port_count[1613],env.pf_vf_mux_scbd_1613.packet_count,1613);
      packet_count_check(port_count[1614],env.pf_vf_mux_scbd_1614.packet_count,1614);
      packet_count_check(port_count[1615],env.pf_vf_mux_scbd_1615.packet_count,1615);
      packet_count_check(port_count[1616],env.pf_vf_mux_scbd_1616.packet_count,1616);
      packet_count_check(port_count[1617],env.pf_vf_mux_scbd_1617.packet_count,1617);
      packet_count_check(port_count[1618],env.pf_vf_mux_scbd_1618.packet_count,1618);
      packet_count_check(port_count[1619],env.pf_vf_mux_scbd_1619.packet_count,1619);
      packet_count_check(port_count[1620],env.pf_vf_mux_scbd_1620.packet_count,1620);
      packet_count_check(port_count[1621],env.pf_vf_mux_scbd_1621.packet_count,1621);
      packet_count_check(port_count[1622],env.pf_vf_mux_scbd_1622.packet_count,1622);
      packet_count_check(port_count[1623],env.pf_vf_mux_scbd_1623.packet_count,1623);
      packet_count_check(port_count[1624],env.pf_vf_mux_scbd_1624.packet_count,1624);
      packet_count_check(port_count[1625],env.pf_vf_mux_scbd_1625.packet_count,1625);
      packet_count_check(port_count[1626],env.pf_vf_mux_scbd_1626.packet_count,1626);
      packet_count_check(port_count[1627],env.pf_vf_mux_scbd_1627.packet_count,1627);
      packet_count_check(port_count[1628],env.pf_vf_mux_scbd_1628.packet_count,1628);
      packet_count_check(port_count[1629],env.pf_vf_mux_scbd_1629.packet_count,1629);
      packet_count_check(port_count[1630],env.pf_vf_mux_scbd_1630.packet_count,1630);
      packet_count_check(port_count[1631],env.pf_vf_mux_scbd_1631.packet_count,1631);
      packet_count_check(port_count[1632],env.pf_vf_mux_scbd_1632.packet_count,1632);
      packet_count_check(port_count[1633],env.pf_vf_mux_scbd_1633.packet_count,1633);
      packet_count_check(port_count[1634],env.pf_vf_mux_scbd_1634.packet_count,1634);
      packet_count_check(port_count[1635],env.pf_vf_mux_scbd_1635.packet_count,1635);
      packet_count_check(port_count[1636],env.pf_vf_mux_scbd_1636.packet_count,1636);
      packet_count_check(port_count[1637],env.pf_vf_mux_scbd_1637.packet_count,1637);
      packet_count_check(port_count[1638],env.pf_vf_mux_scbd_1638.packet_count,1638);
      packet_count_check(port_count[1639],env.pf_vf_mux_scbd_1639.packet_count,1639);
      packet_count_check(port_count[1640],env.pf_vf_mux_scbd_1640.packet_count,1640);
      packet_count_check(port_count[1641],env.pf_vf_mux_scbd_1641.packet_count,1641);
      packet_count_check(port_count[1642],env.pf_vf_mux_scbd_1642.packet_count,1642);
      packet_count_check(port_count[1643],env.pf_vf_mux_scbd_1643.packet_count,1643);
      packet_count_check(port_count[1644],env.pf_vf_mux_scbd_1644.packet_count,1644);
      packet_count_check(port_count[1645],env.pf_vf_mux_scbd_1645.packet_count,1645);
      packet_count_check(port_count[1646],env.pf_vf_mux_scbd_1646.packet_count,1646);
      packet_count_check(port_count[1647],env.pf_vf_mux_scbd_1647.packet_count,1647);
      packet_count_check(port_count[1648],env.pf_vf_mux_scbd_1648.packet_count,1648);
      packet_count_check(port_count[1649],env.pf_vf_mux_scbd_1649.packet_count,1649);
      packet_count_check(port_count[1650],env.pf_vf_mux_scbd_1650.packet_count,1650);
      packet_count_check(port_count[1651],env.pf_vf_mux_scbd_1651.packet_count,1651);
      packet_count_check(port_count[1652],env.pf_vf_mux_scbd_1652.packet_count,1652);
      packet_count_check(port_count[1653],env.pf_vf_mux_scbd_1653.packet_count,1653);
      packet_count_check(port_count[1654],env.pf_vf_mux_scbd_1654.packet_count,1654);
      packet_count_check(port_count[1655],env.pf_vf_mux_scbd_1655.packet_count,1655);
      packet_count_check(port_count[1656],env.pf_vf_mux_scbd_1656.packet_count,1656);
      packet_count_check(port_count[1657],env.pf_vf_mux_scbd_1657.packet_count,1657);
      packet_count_check(port_count[1658],env.pf_vf_mux_scbd_1658.packet_count,1658);
      packet_count_check(port_count[1659],env.pf_vf_mux_scbd_1659.packet_count,1659);
      packet_count_check(port_count[1660],env.pf_vf_mux_scbd_1660.packet_count,1660);
      packet_count_check(port_count[1661],env.pf_vf_mux_scbd_1661.packet_count,1661);
      packet_count_check(port_count[1662],env.pf_vf_mux_scbd_1662.packet_count,1662);
      packet_count_check(port_count[1663],env.pf_vf_mux_scbd_1663.packet_count,1663);
      packet_count_check(port_count[1664],env.pf_vf_mux_scbd_1664.packet_count,1664);
      packet_count_check(port_count[1665],env.pf_vf_mux_scbd_1665.packet_count,1665);
      packet_count_check(port_count[1666],env.pf_vf_mux_scbd_1666.packet_count,1666);
      packet_count_check(port_count[1667],env.pf_vf_mux_scbd_1667.packet_count,1667);
      packet_count_check(port_count[1668],env.pf_vf_mux_scbd_1668.packet_count,1668);
      packet_count_check(port_count[1669],env.pf_vf_mux_scbd_1669.packet_count,1669);
      packet_count_check(port_count[1670],env.pf_vf_mux_scbd_1670.packet_count,1670);
      packet_count_check(port_count[1671],env.pf_vf_mux_scbd_1671.packet_count,1671);
      packet_count_check(port_count[1672],env.pf_vf_mux_scbd_1672.packet_count,1672);
      packet_count_check(port_count[1673],env.pf_vf_mux_scbd_1673.packet_count,1673);
      packet_count_check(port_count[1674],env.pf_vf_mux_scbd_1674.packet_count,1674);
      packet_count_check(port_count[1675],env.pf_vf_mux_scbd_1675.packet_count,1675);
      packet_count_check(port_count[1676],env.pf_vf_mux_scbd_1676.packet_count,1676);
      packet_count_check(port_count[1677],env.pf_vf_mux_scbd_1677.packet_count,1677);
      packet_count_check(port_count[1678],env.pf_vf_mux_scbd_1678.packet_count,1678);
      packet_count_check(port_count[1679],env.pf_vf_mux_scbd_1679.packet_count,1679);
      packet_count_check(port_count[1680],env.pf_vf_mux_scbd_1680.packet_count,1680);
      packet_count_check(port_count[1681],env.pf_vf_mux_scbd_1681.packet_count,1681);
      packet_count_check(port_count[1682],env.pf_vf_mux_scbd_1682.packet_count,1682);
      packet_count_check(port_count[1683],env.pf_vf_mux_scbd_1683.packet_count,1683);
      packet_count_check(port_count[1684],env.pf_vf_mux_scbd_1684.packet_count,1684);
      packet_count_check(port_count[1685],env.pf_vf_mux_scbd_1685.packet_count,1685);
      packet_count_check(port_count[1686],env.pf_vf_mux_scbd_1686.packet_count,1686);
      packet_count_check(port_count[1687],env.pf_vf_mux_scbd_1687.packet_count,1687);
      packet_count_check(port_count[1688],env.pf_vf_mux_scbd_1688.packet_count,1688);
      packet_count_check(port_count[1689],env.pf_vf_mux_scbd_1689.packet_count,1689);
      packet_count_check(port_count[1690],env.pf_vf_mux_scbd_1690.packet_count,1690);
      packet_count_check(port_count[1691],env.pf_vf_mux_scbd_1691.packet_count,1691);
      packet_count_check(port_count[1692],env.pf_vf_mux_scbd_1692.packet_count,1692);
      packet_count_check(port_count[1693],env.pf_vf_mux_scbd_1693.packet_count,1693);
      packet_count_check(port_count[1694],env.pf_vf_mux_scbd_1694.packet_count,1694);
      packet_count_check(port_count[1695],env.pf_vf_mux_scbd_1695.packet_count,1695);
      packet_count_check(port_count[1696],env.pf_vf_mux_scbd_1696.packet_count,1696);
      packet_count_check(port_count[1697],env.pf_vf_mux_scbd_1697.packet_count,1697);
      packet_count_check(port_count[1698],env.pf_vf_mux_scbd_1698.packet_count,1698);
      packet_count_check(port_count[1699],env.pf_vf_mux_scbd_1699.packet_count,1699);
      packet_count_check(port_count[1700],env.pf_vf_mux_scbd_1700.packet_count,1700);
      packet_count_check(port_count[1701],env.pf_vf_mux_scbd_1701.packet_count,1701);
      packet_count_check(port_count[1702],env.pf_vf_mux_scbd_1702.packet_count,1702);
      packet_count_check(port_count[1703],env.pf_vf_mux_scbd_1703.packet_count,1703);
      packet_count_check(port_count[1704],env.pf_vf_mux_scbd_1704.packet_count,1704);
      packet_count_check(port_count[1705],env.pf_vf_mux_scbd_1705.packet_count,1705);
      packet_count_check(port_count[1706],env.pf_vf_mux_scbd_1706.packet_count,1706);
      packet_count_check(port_count[1707],env.pf_vf_mux_scbd_1707.packet_count,1707);
      packet_count_check(port_count[1708],env.pf_vf_mux_scbd_1708.packet_count,1708);
      packet_count_check(port_count[1709],env.pf_vf_mux_scbd_1709.packet_count,1709);
      packet_count_check(port_count[1710],env.pf_vf_mux_scbd_1710.packet_count,1710);
      packet_count_check(port_count[1711],env.pf_vf_mux_scbd_1711.packet_count,1711);
      packet_count_check(port_count[1712],env.pf_vf_mux_scbd_1712.packet_count,1712);
      packet_count_check(port_count[1713],env.pf_vf_mux_scbd_1713.packet_count,1713);
      packet_count_check(port_count[1714],env.pf_vf_mux_scbd_1714.packet_count,1714);
      packet_count_check(port_count[1715],env.pf_vf_mux_scbd_1715.packet_count,1715);
      packet_count_check(port_count[1716],env.pf_vf_mux_scbd_1716.packet_count,1716);
      packet_count_check(port_count[1717],env.pf_vf_mux_scbd_1717.packet_count,1717);
      packet_count_check(port_count[1718],env.pf_vf_mux_scbd_1718.packet_count,1718);
      packet_count_check(port_count[1719],env.pf_vf_mux_scbd_1719.packet_count,1719);
      packet_count_check(port_count[1720],env.pf_vf_mux_scbd_1720.packet_count,1720);
      packet_count_check(port_count[1721],env.pf_vf_mux_scbd_1721.packet_count,1721);
      packet_count_check(port_count[1722],env.pf_vf_mux_scbd_1722.packet_count,1722);
      packet_count_check(port_count[1723],env.pf_vf_mux_scbd_1723.packet_count,1723);
      packet_count_check(port_count[1724],env.pf_vf_mux_scbd_1724.packet_count,1724);
      packet_count_check(port_count[1725],env.pf_vf_mux_scbd_1725.packet_count,1725);
      packet_count_check(port_count[1726],env.pf_vf_mux_scbd_1726.packet_count,1726);
      packet_count_check(port_count[1727],env.pf_vf_mux_scbd_1727.packet_count,1727);
      packet_count_check(port_count[1728],env.pf_vf_mux_scbd_1728.packet_count,1728);
      packet_count_check(port_count[1729],env.pf_vf_mux_scbd_1729.packet_count,1729);
      packet_count_check(port_count[1730],env.pf_vf_mux_scbd_1730.packet_count,1730);
      packet_count_check(port_count[1731],env.pf_vf_mux_scbd_1731.packet_count,1731);
      packet_count_check(port_count[1732],env.pf_vf_mux_scbd_1732.packet_count,1732);
      packet_count_check(port_count[1733],env.pf_vf_mux_scbd_1733.packet_count,1733);
      packet_count_check(port_count[1734],env.pf_vf_mux_scbd_1734.packet_count,1734);
      packet_count_check(port_count[1735],env.pf_vf_mux_scbd_1735.packet_count,1735);
      packet_count_check(port_count[1736],env.pf_vf_mux_scbd_1736.packet_count,1736);
      packet_count_check(port_count[1737],env.pf_vf_mux_scbd_1737.packet_count,1737);
      packet_count_check(port_count[1738],env.pf_vf_mux_scbd_1738.packet_count,1738);
      packet_count_check(port_count[1739],env.pf_vf_mux_scbd_1739.packet_count,1739);
      packet_count_check(port_count[1740],env.pf_vf_mux_scbd_1740.packet_count,1740);
      packet_count_check(port_count[1741],env.pf_vf_mux_scbd_1741.packet_count,1741);
      packet_count_check(port_count[1742],env.pf_vf_mux_scbd_1742.packet_count,1742);
      packet_count_check(port_count[1743],env.pf_vf_mux_scbd_1743.packet_count,1743);
      packet_count_check(port_count[1744],env.pf_vf_mux_scbd_1744.packet_count,1744);
      packet_count_check(port_count[1745],env.pf_vf_mux_scbd_1745.packet_count,1745);
      packet_count_check(port_count[1746],env.pf_vf_mux_scbd_1746.packet_count,1746);
      packet_count_check(port_count[1747],env.pf_vf_mux_scbd_1747.packet_count,1747);
      packet_count_check(port_count[1748],env.pf_vf_mux_scbd_1748.packet_count,1748);
      packet_count_check(port_count[1749],env.pf_vf_mux_scbd_1749.packet_count,1749);
      packet_count_check(port_count[1750],env.pf_vf_mux_scbd_1750.packet_count,1750);
      packet_count_check(port_count[1751],env.pf_vf_mux_scbd_1751.packet_count,1751);
      packet_count_check(port_count[1752],env.pf_vf_mux_scbd_1752.packet_count,1752);
      packet_count_check(port_count[1753],env.pf_vf_mux_scbd_1753.packet_count,1753);
      packet_count_check(port_count[1754],env.pf_vf_mux_scbd_1754.packet_count,1754);
      packet_count_check(port_count[1755],env.pf_vf_mux_scbd_1755.packet_count,1755);
      packet_count_check(port_count[1756],env.pf_vf_mux_scbd_1756.packet_count,1756);
      packet_count_check(port_count[1757],env.pf_vf_mux_scbd_1757.packet_count,1757);
      packet_count_check(port_count[1758],env.pf_vf_mux_scbd_1758.packet_count,1758);
      packet_count_check(port_count[1759],env.pf_vf_mux_scbd_1759.packet_count,1759);
      packet_count_check(port_count[1760],env.pf_vf_mux_scbd_1760.packet_count,1760);
      packet_count_check(port_count[1761],env.pf_vf_mux_scbd_1761.packet_count,1761);
      packet_count_check(port_count[1762],env.pf_vf_mux_scbd_1762.packet_count,1762);
      packet_count_check(port_count[1763],env.pf_vf_mux_scbd_1763.packet_count,1763);
      packet_count_check(port_count[1764],env.pf_vf_mux_scbd_1764.packet_count,1764);
      packet_count_check(port_count[1765],env.pf_vf_mux_scbd_1765.packet_count,1765);
      packet_count_check(port_count[1766],env.pf_vf_mux_scbd_1766.packet_count,1766);
      packet_count_check(port_count[1767],env.pf_vf_mux_scbd_1767.packet_count,1767);
      packet_count_check(port_count[1768],env.pf_vf_mux_scbd_1768.packet_count,1768);
      packet_count_check(port_count[1769],env.pf_vf_mux_scbd_1769.packet_count,1769);
      packet_count_check(port_count[1770],env.pf_vf_mux_scbd_1770.packet_count,1770);
      packet_count_check(port_count[1771],env.pf_vf_mux_scbd_1771.packet_count,1771);
      packet_count_check(port_count[1772],env.pf_vf_mux_scbd_1772.packet_count,1772);
      packet_count_check(port_count[1773],env.pf_vf_mux_scbd_1773.packet_count,1773);
      packet_count_check(port_count[1774],env.pf_vf_mux_scbd_1774.packet_count,1774);
      packet_count_check(port_count[1775],env.pf_vf_mux_scbd_1775.packet_count,1775);
      packet_count_check(port_count[1776],env.pf_vf_mux_scbd_1776.packet_count,1776);
      packet_count_check(port_count[1777],env.pf_vf_mux_scbd_1777.packet_count,1777);
      packet_count_check(port_count[1778],env.pf_vf_mux_scbd_1778.packet_count,1778);
      packet_count_check(port_count[1779],env.pf_vf_mux_scbd_1779.packet_count,1779);
      packet_count_check(port_count[1780],env.pf_vf_mux_scbd_1780.packet_count,1780);
      packet_count_check(port_count[1781],env.pf_vf_mux_scbd_1781.packet_count,1781);
      packet_count_check(port_count[1782],env.pf_vf_mux_scbd_1782.packet_count,1782);
      packet_count_check(port_count[1783],env.pf_vf_mux_scbd_1783.packet_count,1783);
      packet_count_check(port_count[1784],env.pf_vf_mux_scbd_1784.packet_count,1784);
      packet_count_check(port_count[1785],env.pf_vf_mux_scbd_1785.packet_count,1785);
      packet_count_check(port_count[1786],env.pf_vf_mux_scbd_1786.packet_count,1786);
      packet_count_check(port_count[1787],env.pf_vf_mux_scbd_1787.packet_count,1787);
      packet_count_check(port_count[1788],env.pf_vf_mux_scbd_1788.packet_count,1788);
      packet_count_check(port_count[1789],env.pf_vf_mux_scbd_1789.packet_count,1789);
      packet_count_check(port_count[1790],env.pf_vf_mux_scbd_1790.packet_count,1790);
      packet_count_check(port_count[1791],env.pf_vf_mux_scbd_1791.packet_count,1791);
      packet_count_check(port_count[1792],env.pf_vf_mux_scbd_1792.packet_count,1792);
      packet_count_check(port_count[1793],env.pf_vf_mux_scbd_1793.packet_count,1793);
      packet_count_check(port_count[1794],env.pf_vf_mux_scbd_1794.packet_count,1794);
      packet_count_check(port_count[1795],env.pf_vf_mux_scbd_1795.packet_count,1795);
      packet_count_check(port_count[1796],env.pf_vf_mux_scbd_1796.packet_count,1796);
      packet_count_check(port_count[1797],env.pf_vf_mux_scbd_1797.packet_count,1797);
      packet_count_check(port_count[1798],env.pf_vf_mux_scbd_1798.packet_count,1798);
      packet_count_check(port_count[1799],env.pf_vf_mux_scbd_1799.packet_count,1799);
      packet_count_check(port_count[1800],env.pf_vf_mux_scbd_1800.packet_count,1800);
      packet_count_check(port_count[1801],env.pf_vf_mux_scbd_1801.packet_count,1801);
      packet_count_check(port_count[1802],env.pf_vf_mux_scbd_1802.packet_count,1802);
      packet_count_check(port_count[1803],env.pf_vf_mux_scbd_1803.packet_count,1803);
      packet_count_check(port_count[1804],env.pf_vf_mux_scbd_1804.packet_count,1804);
      packet_count_check(port_count[1805],env.pf_vf_mux_scbd_1805.packet_count,1805);
      packet_count_check(port_count[1806],env.pf_vf_mux_scbd_1806.packet_count,1806);
      packet_count_check(port_count[1807],env.pf_vf_mux_scbd_1807.packet_count,1807);
      packet_count_check(port_count[1808],env.pf_vf_mux_scbd_1808.packet_count,1808);
      packet_count_check(port_count[1809],env.pf_vf_mux_scbd_1809.packet_count,1809);
      packet_count_check(port_count[1810],env.pf_vf_mux_scbd_1810.packet_count,1810);
      packet_count_check(port_count[1811],env.pf_vf_mux_scbd_1811.packet_count,1811);
      packet_count_check(port_count[1812],env.pf_vf_mux_scbd_1812.packet_count,1812);
      packet_count_check(port_count[1813],env.pf_vf_mux_scbd_1813.packet_count,1813);
      packet_count_check(port_count[1814],env.pf_vf_mux_scbd_1814.packet_count,1814);
      packet_count_check(port_count[1815],env.pf_vf_mux_scbd_1815.packet_count,1815);
      packet_count_check(port_count[1816],env.pf_vf_mux_scbd_1816.packet_count,1816);
      packet_count_check(port_count[1817],env.pf_vf_mux_scbd_1817.packet_count,1817);
      packet_count_check(port_count[1818],env.pf_vf_mux_scbd_1818.packet_count,1818);
      packet_count_check(port_count[1819],env.pf_vf_mux_scbd_1819.packet_count,1819);
      packet_count_check(port_count[1820],env.pf_vf_mux_scbd_1820.packet_count,1820);
      packet_count_check(port_count[1821],env.pf_vf_mux_scbd_1821.packet_count,1821);
      packet_count_check(port_count[1822],env.pf_vf_mux_scbd_1822.packet_count,1822);
      packet_count_check(port_count[1823],env.pf_vf_mux_scbd_1823.packet_count,1823);
      packet_count_check(port_count[1824],env.pf_vf_mux_scbd_1824.packet_count,1824);
      packet_count_check(port_count[1825],env.pf_vf_mux_scbd_1825.packet_count,1825);
      packet_count_check(port_count[1826],env.pf_vf_mux_scbd_1826.packet_count,1826);
      packet_count_check(port_count[1827],env.pf_vf_mux_scbd_1827.packet_count,1827);
      packet_count_check(port_count[1828],env.pf_vf_mux_scbd_1828.packet_count,1828);
      packet_count_check(port_count[1829],env.pf_vf_mux_scbd_1829.packet_count,1829);
      packet_count_check(port_count[1830],env.pf_vf_mux_scbd_1830.packet_count,1830);
      packet_count_check(port_count[1831],env.pf_vf_mux_scbd_1831.packet_count,1831);
      packet_count_check(port_count[1832],env.pf_vf_mux_scbd_1832.packet_count,1832);
      packet_count_check(port_count[1833],env.pf_vf_mux_scbd_1833.packet_count,1833);
      packet_count_check(port_count[1834],env.pf_vf_mux_scbd_1834.packet_count,1834);
      packet_count_check(port_count[1835],env.pf_vf_mux_scbd_1835.packet_count,1835);
      packet_count_check(port_count[1836],env.pf_vf_mux_scbd_1836.packet_count,1836);
      packet_count_check(port_count[1837],env.pf_vf_mux_scbd_1837.packet_count,1837);
      packet_count_check(port_count[1838],env.pf_vf_mux_scbd_1838.packet_count,1838);
      packet_count_check(port_count[1839],env.pf_vf_mux_scbd_1839.packet_count,1839);
      packet_count_check(port_count[1840],env.pf_vf_mux_scbd_1840.packet_count,1840);
      packet_count_check(port_count[1841],env.pf_vf_mux_scbd_1841.packet_count,1841);
      packet_count_check(port_count[1842],env.pf_vf_mux_scbd_1842.packet_count,1842);
      packet_count_check(port_count[1843],env.pf_vf_mux_scbd_1843.packet_count,1843);
      packet_count_check(port_count[1844],env.pf_vf_mux_scbd_1844.packet_count,1844);
      packet_count_check(port_count[1845],env.pf_vf_mux_scbd_1845.packet_count,1845);
      packet_count_check(port_count[1846],env.pf_vf_mux_scbd_1846.packet_count,1846);
      packet_count_check(port_count[1847],env.pf_vf_mux_scbd_1847.packet_count,1847);
      packet_count_check(port_count[1848],env.pf_vf_mux_scbd_1848.packet_count,1848);
      packet_count_check(port_count[1849],env.pf_vf_mux_scbd_1849.packet_count,1849);
      packet_count_check(port_count[1850],env.pf_vf_mux_scbd_1850.packet_count,1850);
      packet_count_check(port_count[1851],env.pf_vf_mux_scbd_1851.packet_count,1851);
      packet_count_check(port_count[1852],env.pf_vf_mux_scbd_1852.packet_count,1852);
      packet_count_check(port_count[1853],env.pf_vf_mux_scbd_1853.packet_count,1853);
      packet_count_check(port_count[1854],env.pf_vf_mux_scbd_1854.packet_count,1854);
      packet_count_check(port_count[1855],env.pf_vf_mux_scbd_1855.packet_count,1855);
      packet_count_check(port_count[1856],env.pf_vf_mux_scbd_1856.packet_count,1856);
      packet_count_check(port_count[1857],env.pf_vf_mux_scbd_1857.packet_count,1857);
      packet_count_check(port_count[1858],env.pf_vf_mux_scbd_1858.packet_count,1858);
      packet_count_check(port_count[1859],env.pf_vf_mux_scbd_1859.packet_count,1859);
      packet_count_check(port_count[1860],env.pf_vf_mux_scbd_1860.packet_count,1860);
      packet_count_check(port_count[1861],env.pf_vf_mux_scbd_1861.packet_count,1861);
      packet_count_check(port_count[1862],env.pf_vf_mux_scbd_1862.packet_count,1862);
      packet_count_check(port_count[1863],env.pf_vf_mux_scbd_1863.packet_count,1863);
      packet_count_check(port_count[1864],env.pf_vf_mux_scbd_1864.packet_count,1864);
      packet_count_check(port_count[1865],env.pf_vf_mux_scbd_1865.packet_count,1865);
      packet_count_check(port_count[1866],env.pf_vf_mux_scbd_1866.packet_count,1866);
      packet_count_check(port_count[1867],env.pf_vf_mux_scbd_1867.packet_count,1867);
      packet_count_check(port_count[1868],env.pf_vf_mux_scbd_1868.packet_count,1868);
      packet_count_check(port_count[1869],env.pf_vf_mux_scbd_1869.packet_count,1869);
      packet_count_check(port_count[1870],env.pf_vf_mux_scbd_1870.packet_count,1870);
      packet_count_check(port_count[1871],env.pf_vf_mux_scbd_1871.packet_count,1871);
      packet_count_check(port_count[1872],env.pf_vf_mux_scbd_1872.packet_count,1872);
      packet_count_check(port_count[1873],env.pf_vf_mux_scbd_1873.packet_count,1873);
      packet_count_check(port_count[1874],env.pf_vf_mux_scbd_1874.packet_count,1874);
      packet_count_check(port_count[1875],env.pf_vf_mux_scbd_1875.packet_count,1875);
      packet_count_check(port_count[1876],env.pf_vf_mux_scbd_1876.packet_count,1876);
      packet_count_check(port_count[1877],env.pf_vf_mux_scbd_1877.packet_count,1877);
      packet_count_check(port_count[1878],env.pf_vf_mux_scbd_1878.packet_count,1878);
      packet_count_check(port_count[1879],env.pf_vf_mux_scbd_1879.packet_count,1879);
      packet_count_check(port_count[1880],env.pf_vf_mux_scbd_1880.packet_count,1880);
      packet_count_check(port_count[1881],env.pf_vf_mux_scbd_1881.packet_count,1881);
      packet_count_check(port_count[1882],env.pf_vf_mux_scbd_1882.packet_count,1882);
      packet_count_check(port_count[1883],env.pf_vf_mux_scbd_1883.packet_count,1883);
      packet_count_check(port_count[1884],env.pf_vf_mux_scbd_1884.packet_count,1884);
      packet_count_check(port_count[1885],env.pf_vf_mux_scbd_1885.packet_count,1885);
      packet_count_check(port_count[1886],env.pf_vf_mux_scbd_1886.packet_count,1886);
      packet_count_check(port_count[1887],env.pf_vf_mux_scbd_1887.packet_count,1887);
      packet_count_check(port_count[1888],env.pf_vf_mux_scbd_1888.packet_count,1888);
      packet_count_check(port_count[1889],env.pf_vf_mux_scbd_1889.packet_count,1889);
      packet_count_check(port_count[1890],env.pf_vf_mux_scbd_1890.packet_count,1890);
      packet_count_check(port_count[1891],env.pf_vf_mux_scbd_1891.packet_count,1891);
      packet_count_check(port_count[1892],env.pf_vf_mux_scbd_1892.packet_count,1892);
      packet_count_check(port_count[1893],env.pf_vf_mux_scbd_1893.packet_count,1893);
      packet_count_check(port_count[1894],env.pf_vf_mux_scbd_1894.packet_count,1894);
      packet_count_check(port_count[1895],env.pf_vf_mux_scbd_1895.packet_count,1895);
      packet_count_check(port_count[1896],env.pf_vf_mux_scbd_1896.packet_count,1896);
      packet_count_check(port_count[1897],env.pf_vf_mux_scbd_1897.packet_count,1897);
      packet_count_check(port_count[1898],env.pf_vf_mux_scbd_1898.packet_count,1898);
      packet_count_check(port_count[1899],env.pf_vf_mux_scbd_1899.packet_count,1899);
      packet_count_check(port_count[1900],env.pf_vf_mux_scbd_1900.packet_count,1900);
      packet_count_check(port_count[1901],env.pf_vf_mux_scbd_1901.packet_count,1901);
      packet_count_check(port_count[1902],env.pf_vf_mux_scbd_1902.packet_count,1902);
      packet_count_check(port_count[1903],env.pf_vf_mux_scbd_1903.packet_count,1903);
      packet_count_check(port_count[1904],env.pf_vf_mux_scbd_1904.packet_count,1904);
      packet_count_check(port_count[1905],env.pf_vf_mux_scbd_1905.packet_count,1905);
      packet_count_check(port_count[1906],env.pf_vf_mux_scbd_1906.packet_count,1906);
      packet_count_check(port_count[1907],env.pf_vf_mux_scbd_1907.packet_count,1907);
      packet_count_check(port_count[1908],env.pf_vf_mux_scbd_1908.packet_count,1908);
      packet_count_check(port_count[1909],env.pf_vf_mux_scbd_1909.packet_count,1909);
      packet_count_check(port_count[1910],env.pf_vf_mux_scbd_1910.packet_count,1910);
      packet_count_check(port_count[1911],env.pf_vf_mux_scbd_1911.packet_count,1911);
      packet_count_check(port_count[1912],env.pf_vf_mux_scbd_1912.packet_count,1912);
      packet_count_check(port_count[1913],env.pf_vf_mux_scbd_1913.packet_count,1913);
      packet_count_check(port_count[1914],env.pf_vf_mux_scbd_1914.packet_count,1914);
      packet_count_check(port_count[1915],env.pf_vf_mux_scbd_1915.packet_count,1915);
      packet_count_check(port_count[1916],env.pf_vf_mux_scbd_1916.packet_count,1916);
      packet_count_check(port_count[1917],env.pf_vf_mux_scbd_1917.packet_count,1917);
      packet_count_check(port_count[1918],env.pf_vf_mux_scbd_1918.packet_count,1918);
      packet_count_check(port_count[1919],env.pf_vf_mux_scbd_1919.packet_count,1919);
      packet_count_check(port_count[1920],env.pf_vf_mux_scbd_1920.packet_count,1920);
      packet_count_check(port_count[1921],env.pf_vf_mux_scbd_1921.packet_count,1921);
      packet_count_check(port_count[1922],env.pf_vf_mux_scbd_1922.packet_count,1922);
      packet_count_check(port_count[1923],env.pf_vf_mux_scbd_1923.packet_count,1923);
      packet_count_check(port_count[1924],env.pf_vf_mux_scbd_1924.packet_count,1924);
      packet_count_check(port_count[1925],env.pf_vf_mux_scbd_1925.packet_count,1925);
      packet_count_check(port_count[1926],env.pf_vf_mux_scbd_1926.packet_count,1926);
      packet_count_check(port_count[1927],env.pf_vf_mux_scbd_1927.packet_count,1927);
      packet_count_check(port_count[1928],env.pf_vf_mux_scbd_1928.packet_count,1928);
      packet_count_check(port_count[1929],env.pf_vf_mux_scbd_1929.packet_count,1929);
      packet_count_check(port_count[1930],env.pf_vf_mux_scbd_1930.packet_count,1930);
      packet_count_check(port_count[1931],env.pf_vf_mux_scbd_1931.packet_count,1931);
      packet_count_check(port_count[1932],env.pf_vf_mux_scbd_1932.packet_count,1932);
      packet_count_check(port_count[1933],env.pf_vf_mux_scbd_1933.packet_count,1933);
      packet_count_check(port_count[1934],env.pf_vf_mux_scbd_1934.packet_count,1934);
      packet_count_check(port_count[1935],env.pf_vf_mux_scbd_1935.packet_count,1935);
      packet_count_check(port_count[1936],env.pf_vf_mux_scbd_1936.packet_count,1936);
      packet_count_check(port_count[1937],env.pf_vf_mux_scbd_1937.packet_count,1937);
      packet_count_check(port_count[1938],env.pf_vf_mux_scbd_1938.packet_count,1938);
      packet_count_check(port_count[1939],env.pf_vf_mux_scbd_1939.packet_count,1939);
      packet_count_check(port_count[1940],env.pf_vf_mux_scbd_1940.packet_count,1940);
      packet_count_check(port_count[1941],env.pf_vf_mux_scbd_1941.packet_count,1941);
      packet_count_check(port_count[1942],env.pf_vf_mux_scbd_1942.packet_count,1942);
      packet_count_check(port_count[1943],env.pf_vf_mux_scbd_1943.packet_count,1943);
      packet_count_check(port_count[1944],env.pf_vf_mux_scbd_1944.packet_count,1944);
      packet_count_check(port_count[1945],env.pf_vf_mux_scbd_1945.packet_count,1945);
      packet_count_check(port_count[1946],env.pf_vf_mux_scbd_1946.packet_count,1946);
      packet_count_check(port_count[1947],env.pf_vf_mux_scbd_1947.packet_count,1947);
      packet_count_check(port_count[1948],env.pf_vf_mux_scbd_1948.packet_count,1948);
      packet_count_check(port_count[1949],env.pf_vf_mux_scbd_1949.packet_count,1949);
      packet_count_check(port_count[1950],env.pf_vf_mux_scbd_1950.packet_count,1950);
      packet_count_check(port_count[1951],env.pf_vf_mux_scbd_1951.packet_count,1951);
      packet_count_check(port_count[1952],env.pf_vf_mux_scbd_1952.packet_count,1952);
      packet_count_check(port_count[1953],env.pf_vf_mux_scbd_1953.packet_count,1953);
      packet_count_check(port_count[1954],env.pf_vf_mux_scbd_1954.packet_count,1954);
      packet_count_check(port_count[1955],env.pf_vf_mux_scbd_1955.packet_count,1955);
      packet_count_check(port_count[1956],env.pf_vf_mux_scbd_1956.packet_count,1956);
      packet_count_check(port_count[1957],env.pf_vf_mux_scbd_1957.packet_count,1957);
      packet_count_check(port_count[1958],env.pf_vf_mux_scbd_1958.packet_count,1958);
      packet_count_check(port_count[1959],env.pf_vf_mux_scbd_1959.packet_count,1959);
      packet_count_check(port_count[1960],env.pf_vf_mux_scbd_1960.packet_count,1960);
      packet_count_check(port_count[1961],env.pf_vf_mux_scbd_1961.packet_count,1961);
      packet_count_check(port_count[1962],env.pf_vf_mux_scbd_1962.packet_count,1962);
      packet_count_check(port_count[1963],env.pf_vf_mux_scbd_1963.packet_count,1963);
      packet_count_check(port_count[1964],env.pf_vf_mux_scbd_1964.packet_count,1964);
      packet_count_check(port_count[1965],env.pf_vf_mux_scbd_1965.packet_count,1965);
      packet_count_check(port_count[1966],env.pf_vf_mux_scbd_1966.packet_count,1966);
      packet_count_check(port_count[1967],env.pf_vf_mux_scbd_1967.packet_count,1967);
      packet_count_check(port_count[1968],env.pf_vf_mux_scbd_1968.packet_count,1968);
      packet_count_check(port_count[1969],env.pf_vf_mux_scbd_1969.packet_count,1969);
      packet_count_check(port_count[1970],env.pf_vf_mux_scbd_1970.packet_count,1970);
      packet_count_check(port_count[1971],env.pf_vf_mux_scbd_1971.packet_count,1971);
      packet_count_check(port_count[1972],env.pf_vf_mux_scbd_1972.packet_count,1972);
      packet_count_check(port_count[1973],env.pf_vf_mux_scbd_1973.packet_count,1973);
      packet_count_check(port_count[1974],env.pf_vf_mux_scbd_1974.packet_count,1974);
      packet_count_check(port_count[1975],env.pf_vf_mux_scbd_1975.packet_count,1975);
      packet_count_check(port_count[1976],env.pf_vf_mux_scbd_1976.packet_count,1976);
      packet_count_check(port_count[1977],env.pf_vf_mux_scbd_1977.packet_count,1977);
      packet_count_check(port_count[1978],env.pf_vf_mux_scbd_1978.packet_count,1978);
      packet_count_check(port_count[1979],env.pf_vf_mux_scbd_1979.packet_count,1979);
      packet_count_check(port_count[1980],env.pf_vf_mux_scbd_1980.packet_count,1980);
      packet_count_check(port_count[1981],env.pf_vf_mux_scbd_1981.packet_count,1981);
      packet_count_check(port_count[1982],env.pf_vf_mux_scbd_1982.packet_count,1982);
      packet_count_check(port_count[1983],env.pf_vf_mux_scbd_1983.packet_count,1983);
      packet_count_check(port_count[1984],env.pf_vf_mux_scbd_1984.packet_count,1984);
      packet_count_check(port_count[1985],env.pf_vf_mux_scbd_1985.packet_count,1985);
      packet_count_check(port_count[1986],env.pf_vf_mux_scbd_1986.packet_count,1986);
      packet_count_check(port_count[1987],env.pf_vf_mux_scbd_1987.packet_count,1987);
      packet_count_check(port_count[1988],env.pf_vf_mux_scbd_1988.packet_count,1988);
      packet_count_check(port_count[1989],env.pf_vf_mux_scbd_1989.packet_count,1989);
      packet_count_check(port_count[1990],env.pf_vf_mux_scbd_1990.packet_count,1990);
      packet_count_check(port_count[1991],env.pf_vf_mux_scbd_1991.packet_count,1991);
      packet_count_check(port_count[1992],env.pf_vf_mux_scbd_1992.packet_count,1992);
      packet_count_check(port_count[1993],env.pf_vf_mux_scbd_1993.packet_count,1993);
      packet_count_check(port_count[1994],env.pf_vf_mux_scbd_1994.packet_count,1994);
      packet_count_check(port_count[1995],env.pf_vf_mux_scbd_1995.packet_count,1995);
      packet_count_check(port_count[1996],env.pf_vf_mux_scbd_1996.packet_count,1996);
      packet_count_check(port_count[1997],env.pf_vf_mux_scbd_1997.packet_count,1997);
      packet_count_check(port_count[1998],env.pf_vf_mux_scbd_1998.packet_count,1998);
      packet_count_check(port_count[1999],env.pf_vf_mux_scbd_1999.packet_count,1999);
      packet_count_check(port_count[2000],env.pf_vf_mux_scbd_2000.packet_count,2000);
      packet_count_check(port_count[2001],env.pf_vf_mux_scbd_2001.packet_count,2001);
      packet_count_check(port_count[2002],env.pf_vf_mux_scbd_2002.packet_count,2002);
      packet_count_check(port_count[2003],env.pf_vf_mux_scbd_2003.packet_count,2003);
      packet_count_check(port_count[2004],env.pf_vf_mux_scbd_2004.packet_count,2004);
      packet_count_check(port_count[2005],env.pf_vf_mux_scbd_2005.packet_count,2005);
      packet_count_check(port_count[2006],env.pf_vf_mux_scbd_2006.packet_count,2006);
      packet_count_check(port_count[2007],env.pf_vf_mux_scbd_2007.packet_count,2007);
      packet_count_check(port_count[2008],env.pf_vf_mux_scbd_2008.packet_count,2008);
      packet_count_check(port_count[2009],env.pf_vf_mux_scbd_2009.packet_count,2009);
      packet_count_check(port_count[2010],env.pf_vf_mux_scbd_2010.packet_count,2010);
      packet_count_check(port_count[2011],env.pf_vf_mux_scbd_2011.packet_count,2011);
      packet_count_check(port_count[2012],env.pf_vf_mux_scbd_2012.packet_count,2012);
      packet_count_check(port_count[2013],env.pf_vf_mux_scbd_2013.packet_count,2013);
      packet_count_check(port_count[2014],env.pf_vf_mux_scbd_2014.packet_count,2014);
      packet_count_check(port_count[2015],env.pf_vf_mux_scbd_2015.packet_count,2015);
      packet_count_check(port_count[2016],env.pf_vf_mux_scbd_2016.packet_count,2016);
      packet_count_check(port_count[2017],env.pf_vf_mux_scbd_2017.packet_count,2017);
      packet_count_check(port_count[2018],env.pf_vf_mux_scbd_2018.packet_count,2018);
      packet_count_check(port_count[2019],env.pf_vf_mux_scbd_2019.packet_count,2019);
      packet_count_check(port_count[2020],env.pf_vf_mux_scbd_2020.packet_count,2020);
      packet_count_check(port_count[2021],env.pf_vf_mux_scbd_2021.packet_count,2021);
      packet_count_check(port_count[2022],env.pf_vf_mux_scbd_2022.packet_count,2022);
      packet_count_check(port_count[2023],env.pf_vf_mux_scbd_2023.packet_count,2023);
      packet_count_check(port_count[2024],env.pf_vf_mux_scbd_2024.packet_count,2024);
      packet_count_check(port_count[2025],env.pf_vf_mux_scbd_2025.packet_count,2025);
      packet_count_check(port_count[2026],env.pf_vf_mux_scbd_2026.packet_count,2026);
      packet_count_check(port_count[2027],env.pf_vf_mux_scbd_2027.packet_count,2027);
      packet_count_check(port_count[2028],env.pf_vf_mux_scbd_2028.packet_count,2028);
      packet_count_check(port_count[2029],env.pf_vf_mux_scbd_2029.packet_count,2029);
      packet_count_check(port_count[2030],env.pf_vf_mux_scbd_2030.packet_count,2030);
      packet_count_check(port_count[2031],env.pf_vf_mux_scbd_2031.packet_count,2031);
      packet_count_check(port_count[2032],env.pf_vf_mux_scbd_2032.packet_count,2032);
      packet_count_check(port_count[2033],env.pf_vf_mux_scbd_2033.packet_count,2033);
      packet_count_check(port_count[2034],env.pf_vf_mux_scbd_2034.packet_count,2034);
      packet_count_check(port_count[2035],env.pf_vf_mux_scbd_2035.packet_count,2035);
      packet_count_check(port_count[2036],env.pf_vf_mux_scbd_2036.packet_count,2036);
      packet_count_check(port_count[2037],env.pf_vf_mux_scbd_2037.packet_count,2037);
      packet_count_check(port_count[2038],env.pf_vf_mux_scbd_2038.packet_count,2038);
      packet_count_check(port_count[2039],env.pf_vf_mux_scbd_2039.packet_count,2039);
      packet_count_check(port_count[2040],env.pf_vf_mux_scbd_2040.packet_count,2040);
      packet_count_check(port_count[2041],env.pf_vf_mux_scbd_2041.packet_count,2041);
      packet_count_check(port_count[2042],env.pf_vf_mux_scbd_2042.packet_count,2042);
      packet_count_check(port_count[2043],env.pf_vf_mux_scbd_2043.packet_count,2043);
      packet_count_check(port_count[2044],env.pf_vf_mux_scbd_2044.packet_count,2044);
      packet_count_check(port_count[2045],env.pf_vf_mux_scbd_2045.packet_count,2045);
      packet_count_check(port_count[2046],env.pf_vf_mux_scbd_2046.packet_count,2046);
      packet_count_check(port_count[2047],env.pf_vf_mux_scbd_2047.packet_count,2047);
      `endif
  endfunction

endclass

`endif // GUARD_PF_VF_MUX_BASE_TEST_SV
